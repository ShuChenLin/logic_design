`timescale 1ns/1ps

module Multiplier_4bit(a, b, p);
    input [4-1:0] a, b;
    output [8-1:0] p;

endmodule
