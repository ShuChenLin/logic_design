`timescale 1ns/1ps

module mem_addr_gen(
   input clk,
   input rst,
   input [2:0] state,
   input [9:0] h_cnt,
   input [9:0] v_cnt,
   input [8:0] word_num, // which word to display
   input [5:0] wrong_cnt,
   input [5:0] letter,
   input correct,
   input [10:0] word_cnt, // which word should I type
   input [3:0] cpm1, cpm2, cpm3,
   input cursor,
   output reg [3:0] red, green, blue
   );
   
    parameter WAIT = 3'b000;
    parameter WAIT_TO_START = 3'b001;
    parameter WORD = 3'b010;
    parameter WRONG = 3'b011;
    parameter FINISH = 3'b100;
    
   wire [11:0] Upperletter [1663:0];
   wire [11:0] Lowerletter [1663:0];
   wire [11:0] otherletter [255:0];
   wire [11:0] CPM [13311:0];
   //cpm_digits are for finding the rgb of the number, count_for_cpm is for what to output on the display
   wire [16:0] cpm_digit1, cpm_digit2, cpm_digit3, count_for_cpm, CCPPMM;
   wire [15:0] place, place2, place3;
   
   // variables for find the character in memories====================================================
   assign place = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * letter);
   assign place2 = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * (letter - 26));
   assign place3 = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * (letter - 30));
   assign cpm_digit1 = (h_cnt % 32) + 32 * (v_cnt % 32) + (1024 * (3 + cpm1));
   assign cpm_digit2 = (h_cnt % 32) + 32 * (v_cnt % 32) + (1024 * (3 + cpm2));
   assign cpm_digit3 = (h_cnt % 32) + 32 * (v_cnt % 32) + (1024 * (3 + cpm3));
   assign count_for_cpm = (h_cnt - 224) / 32;
   assign CCPPMM = (count_for_cpm < 3) ? (h_cnt % 32) + 32 * (v_cnt % 32) + (1024 * count_for_cpm) : 0;
   //==================================================================================================
   
   always @(*) begin
        {red, green, blue} = 12'b111111111111;
        if (state == FINISH) begin
            // only CPM in the middle of monitor
            if (v_cnt >= 224 && v_cnt <= 256 && h_cnt >= 224 && h_cnt <= 416) begin
                if (count_for_cpm < 3) begin
                    {red, green, blue} = CPM[CCPPMM];
                end else begin
                    if (count_for_cpm == 5) {red, green, blue} = CPM[cpm_digit1];
                    else if (count_for_cpm == 4) {red, green, blue} = CPM[cpm_digit2];
                    else if (count_for_cpm == 3) {red, green, blue} = CPM[cpm_digit3];
                end
            end
        end
        else begin
            if (h_cnt >= 80 && h_cnt <= 560 && v_cnt >= 208 && v_cnt <= 280) begin
                // place to put the article
                if (word_num > 298 || (v_cnt / 8) == 27 || (v_cnt) / 8 == 29 || (v_cnt) / 8 == 31 || (v_cnt) / 8 == 33 || (v_cnt) / 8 == 35) {red, green, blue} = 12'b111111111111;
                else begin
                    if (correct && (word_num >= word_cnt) && (word_num < word_cnt + wrong_cnt)) begin
                        //wrong words
                        if (letter <= 25) {red, green, blue} = (Lowerletter[place] == 12'b0) ? 12'b0 : 12'b111100110000;
                        else if (letter >= 26 && letter <= 29) {red, green, blue} = (otherletter[place2] == 12'b0) ? 12'b0 : 12'b111100110000;
                        else {red, green, blue} = (Upperletter[place3] == 12'b0) ? 12'b0 : 12'b111100110000;

                    end else if (word_num < word_cnt) begin
                        //already finished words
                        if (letter <= 25) {red, green, blue} = (Lowerletter[place] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;
                        else if (letter >= 26 && letter <= 29) {red, green, blue} = (otherletter[place2] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;
                        else {red, green, blue} = (Upperletter[place3] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;

                    end else begin
                        //word typing, place of cursor
                        if (letter <= 25) {red, green, blue} = (cursor) ? ~Lowerletter[place] : Lowerletter[place];
                        else if (letter >= 26 && letter <= 29) {red, green, blue} = (cursor) ? ~otherletter[place2] : otherletter[place2];
                        else {red, green, blue} = (cursor) ? ~Upperletter[place3] : Upperletter[place3];

                    end
                end
            end else begin
                // output for CPM
                if (v_cnt >= 64 && v_cnt <= 96 && h_cnt >= 224 && h_cnt <= 416) begin
                    if (count_for_cpm < 3) begin
                        {red, green, blue} = CPM[CCPPMM];
                    end else begin
                        if (count_for_cpm == 5) {red, green, blue} = CPM[cpm_digit1];
                        else if (count_for_cpm == 4) {red, green, blue} = CPM[cpm_digit2];
                        else if (count_for_cpm == 3) {red, green, blue} = CPM[cpm_digit3];
                    end
                end
            end
        end
    end


// input the rgb representation of the pictures I want    
assign otherletter[0] = 12'b111111111111;
assign otherletter[1] = 12'b111111111111;
assign otherletter[2] = 12'b111111111111;
assign otherletter[3] = 12'b111111111111;
assign otherletter[4] = 12'b111111111111;
assign otherletter[5] = 12'b111111111111;
assign otherletter[6] = 12'b111111111111;
assign otherletter[7] = 12'b111111111111;
assign otherletter[8] = 12'b111111111111;
assign otherletter[9] = 12'b111111111111;
assign otherletter[10] = 12'b111111111111;
assign otherletter[11] = 12'b111111111111;
assign otherletter[12] = 12'b111111111111;
assign otherletter[13] = 12'b111111111111;
assign otherletter[14] = 12'b111111111111;
assign otherletter[15] = 12'b111111111111;
assign otherletter[16] = 12'b111111111111;
assign otherletter[17] = 12'b111111111111;
assign otherletter[18] = 12'b111111111111;
assign otherletter[19] = 12'b111111111111;
assign otherletter[20] = 12'b111111111111;
assign otherletter[21] = 12'b111111111111;
assign otherletter[22] = 12'b111111111111;
assign otherletter[23] = 12'b111111111111;
assign otherletter[24] = 12'b111111111111;
assign otherletter[25] = 12'b111111111111;
assign otherletter[26] = 12'b111111111111;
assign otherletter[27] = 12'b111111111111;
assign otherletter[28] = 12'b111111111111;
assign otherletter[29] = 12'b111111111111;
assign otherletter[30] = 12'b111111111111;
assign otherletter[31] = 12'b111111111111;
assign otherletter[32] = 12'b111111111111;
assign otherletter[33] = 12'b111111111111;
assign otherletter[34] = 12'b111111111111;
assign otherletter[35] = 12'b111111111111;
assign otherletter[36] = 12'b111111111111;
assign otherletter[37] = 12'b111111111111;
assign otherletter[38] = 12'b111111111111;
assign otherletter[39] = 12'b111111111111;
assign otherletter[40] = 12'b111111111111;
assign otherletter[41] = 12'b111111111111;
assign otherletter[42] = 12'b111111111111;
assign otherletter[43] = 12'b111111111111;
assign otherletter[44] = 12'b111111111111;
assign otherletter[45] = 12'b111111111111;
assign otherletter[46] = 12'b111111111111;
assign otherletter[47] = 12'b111111111111;
assign otherletter[48] = 12'b111111111111;
assign otherletter[49] = 12'b111111111111;
assign otherletter[50] = 12'b111111111111;
assign otherletter[51] = 12'b111111111111;
assign otherletter[52] = 12'b111111111111;
assign otherletter[53] = 12'b111111111111;
assign otherletter[54] = 12'b111111111111;
assign otherletter[55] = 12'b111111111111;
assign otherletter[56] = 12'b111111111111;
assign otherletter[57] = 12'b111111111111;
assign otherletter[58] = 12'b111111111111;
assign otherletter[59] = 12'b111111111111;
assign otherletter[60] = 12'b111111111111;
assign otherletter[61] = 12'b111111111111;
assign otherletter[62] = 12'b111111111111;
assign otherletter[63] = 12'b111111111111;
assign otherletter[64] = 12'b111111111111;
assign otherletter[65] = 12'b111111111111;
assign otherletter[66] = 12'b111111111111;
assign otherletter[67] = 12'b111111111111;
assign otherletter[68] = 12'b111111111111;
assign otherletter[69] = 12'b111111111111;
assign otherletter[70] = 12'b111111111111;
assign otherletter[71] = 12'b111111111111;
assign otherletter[72] = 12'b111111111111;
assign otherletter[73] = 12'b111111111111;
assign otherletter[74] = 12'b111111111111;
assign otherletter[75] = 12'b111111111111;
assign otherletter[76] = 12'b111111111111;
assign otherletter[77] = 12'b111111111111;
assign otherletter[78] = 12'b111111111111;
assign otherletter[79] = 12'b111111111111;
assign otherletter[80] = 12'b111111111111;
assign otherletter[81] = 12'b111111111111;
assign otherletter[82] = 12'b111111111111;
assign otherletter[83] = 12'b111111111111;
assign otherletter[84] = 12'b111111111111;
assign otherletter[85] = 12'b111111111111;
assign otherletter[86] = 12'b111111111111;
assign otherletter[87] = 12'b111111111111;
assign otherletter[88] = 12'b111111111111;
assign otherletter[89] = 12'b111111111111;
assign otherletter[90] = 12'b111111111111;
assign otherletter[91] = 12'b111111111111;
assign otherletter[92] = 12'b111111111111;
assign otherletter[93] = 12'b111111111111;
assign otherletter[94] = 12'b111111111111;
assign otherletter[95] = 12'b111111111111;
assign otherletter[96] = 12'b111111111111;
assign otherletter[97] = 12'b111111111111;
assign otherletter[98] = 12'b111111111111;
assign otherletter[99] = 12'b111111111111;
assign otherletter[100] = 12'b111111111111;
assign otherletter[101] = 12'b111111111111;
assign otherletter[102] = 12'b111111111111;
assign otherletter[103] = 12'b111111111111;
assign otherletter[104] = 12'b111111111111;
assign otherletter[105] = 12'b111111111111;
assign otherletter[106] = 12'b111111111111;
assign otherletter[107] = 12'b111111111111;
assign otherletter[108] = 12'b111111111111;
assign otherletter[109] = 12'b111111111111;
assign otherletter[110] = 12'b111111111111;
assign otherletter[111] = 12'b111111111111;
assign otherletter[112] = 12'b111111111111;
assign otherletter[113] = 12'b111111111111;
assign otherletter[114] = 12'b111111111111;
assign otherletter[115] = 12'b000000000000;
assign otherletter[116] = 12'b111111111111;
assign otherletter[117] = 12'b111111111111;
assign otherletter[118] = 12'b111111111111;
assign otherletter[119] = 12'b111111111111;
assign otherletter[120] = 12'b111111111111;
assign otherletter[121] = 12'b111111111111;
assign otherletter[122] = 12'b111111111111;
assign otherletter[123] = 12'b000000000000;
assign otherletter[124] = 12'b111111111111;
assign otherletter[125] = 12'b111111111111;
assign otherletter[126] = 12'b111111111111;
assign otherletter[127] = 12'b111111111111;
assign otherletter[128] = 12'b111111111111;
assign otherletter[129] = 12'b111111111111;
assign otherletter[130] = 12'b111111111111;
assign otherletter[131] = 12'b111111111111;
assign otherletter[132] = 12'b111111111111;
assign otherletter[133] = 12'b111111111111;
assign otherletter[134] = 12'b111111111111;
assign otherletter[135] = 12'b111111111111;
assign otherletter[136] = 12'b111111111111;
assign otherletter[137] = 12'b111111111111;
assign otherletter[138] = 12'b111111111111;
assign otherletter[139] = 12'b111111111111;
assign otherletter[140] = 12'b111111111111;
assign otherletter[141] = 12'b111111111111;
assign otherletter[142] = 12'b111111111111;
assign otherletter[143] = 12'b111111111111;
assign otherletter[144] = 12'b111111111111;
assign otherletter[145] = 12'b111111111111;
assign otherletter[146] = 12'b111111111111;
assign otherletter[147] = 12'b111111111111;
assign otherletter[148] = 12'b111111111111;
assign otherletter[149] = 12'b111111111111;
assign otherletter[150] = 12'b111111111111;
assign otherletter[151] = 12'b111111111111;
assign otherletter[152] = 12'b111111111111;
assign otherletter[153] = 12'b111111111111;
assign otherletter[154] = 12'b111111111111;
assign otherletter[155] = 12'b111111111111;
assign otherletter[156] = 12'b111111111111;
assign otherletter[157] = 12'b111111111111;
assign otherletter[158] = 12'b111111111111;
assign otherletter[159] = 12'b111111111111;
assign otherletter[160] = 12'b111111111111;
assign otherletter[161] = 12'b111111111111;
assign otherletter[162] = 12'b111111111111;
assign otherletter[163] = 12'b111111111111;
assign otherletter[164] = 12'b111111111111;
assign otherletter[165] = 12'b111111111111;
assign otherletter[166] = 12'b111111111111;
assign otherletter[167] = 12'b111111111111;
assign otherletter[168] = 12'b111111111111;
assign otherletter[169] = 12'b111111111111;
assign otherletter[170] = 12'b111111111111;
assign otherletter[171] = 12'b111111111111;
assign otherletter[172] = 12'b111111111111;
assign otherletter[173] = 12'b111111111111;
assign otherletter[174] = 12'b111111111111;
assign otherletter[175] = 12'b111111111111;
assign otherletter[176] = 12'b111111111111;
assign otherletter[177] = 12'b111111111111;
assign otherletter[178] = 12'b111111111111;
assign otherletter[179] = 12'b000000000000;
assign otherletter[180] = 12'b111111111111;
assign otherletter[181] = 12'b111111111111;
assign otherletter[182] = 12'b111111111111;
assign otherletter[183] = 12'b111111111111;
assign otherletter[184] = 12'b111111111111;
assign otherletter[185] = 12'b111111111111;
assign otherletter[186] = 12'b111111111111;
assign otherletter[187] = 12'b111111111111;
assign otherletter[188] = 12'b111111111111;
assign otherletter[189] = 12'b111111111111;
assign otherletter[190] = 12'b111111111111;
assign otherletter[191] = 12'b111111111111;
assign otherletter[192] = 12'b111111111111;
assign otherletter[193] = 12'b111111111111;
assign otherletter[194] = 12'b111111111111;
assign otherletter[195] = 12'b000000000000;
assign otherletter[196] = 12'b111111111111;
assign otherletter[197] = 12'b111111111111;
assign otherletter[198] = 12'b111111111111;
assign otherletter[199] = 12'b111111111111;
assign otherletter[200] = 12'b111111111111;
assign otherletter[201] = 12'b111111111111;
assign otherletter[202] = 12'b111111111111;
assign otherletter[203] = 12'b000000000000;
assign otherletter[204] = 12'b111111111111;
assign otherletter[205] = 12'b111111111111;
assign otherletter[206] = 12'b111111111111;
assign otherletter[207] = 12'b111111111111;
assign otherletter[208] = 12'b111111111111;
assign otherletter[209] = 12'b111111111111;
assign otherletter[210] = 12'b111111111111;
assign otherletter[211] = 12'b111111111111;
assign otherletter[212] = 12'b111111111111;
assign otherletter[213] = 12'b111111111111;
assign otherletter[214] = 12'b111111111111;
assign otherletter[215] = 12'b111111111111;
assign otherletter[216] = 12'b111111111111;
assign otherletter[217] = 12'b111111111111;
assign otherletter[218] = 12'b111111111111;
assign otherletter[219] = 12'b111111111111;
assign otherletter[220] = 12'b111111111111;
assign otherletter[221] = 12'b111111111111;
assign otherletter[222] = 12'b111111111111;
assign otherletter[223] = 12'b111111111111;
assign otherletter[224] = 12'b111111111111;
assign otherletter[225] = 12'b111111111111;
assign otherletter[226] = 12'b111111111111;
assign otherletter[227] = 12'b111111111111;
assign otherletter[228] = 12'b111111111111;
assign otherletter[229] = 12'b111111111111;
assign otherletter[230] = 12'b111111111111;
assign otherletter[231] = 12'b111111111111;
assign otherletter[232] = 12'b111111111111;
assign otherletter[233] = 12'b111111111111;
assign otherletter[234] = 12'b111111111111;
assign otherletter[235] = 12'b111111111111;
assign otherletter[236] = 12'b111111111111;
assign otherletter[237] = 12'b111111111111;
assign otherletter[238] = 12'b111111111111;
assign otherletter[239] = 12'b111111111111;
assign otherletter[240] = 12'b111111111111;
assign otherletter[241] = 12'b111111111111;
assign otherletter[242] = 12'b111111111111;
assign otherletter[243] = 12'b111111111111;
assign otherletter[244] = 12'b111111111111;
assign otherletter[245] = 12'b111111111111;
assign otherletter[246] = 12'b111111111111;
assign otherletter[247] = 12'b111111111111;
assign otherletter[248] = 12'b111111111111;
assign otherletter[249] = 12'b111111111111;
assign otherletter[250] = 12'b111111111111;
assign otherletter[251] = 12'b111111111111;
assign otherletter[252] = 12'b111111111111;
assign otherletter[253] = 12'b111111111111;
assign otherletter[254] = 12'b111111111111;
assign otherletter[255] = 12'b111111111111;    
assign Lowerletter[0] = 12'b111111111111;
assign Lowerletter[1] = 12'b111111111111;
assign Lowerletter[2] = 12'b111111111111;
assign Lowerletter[3] = 12'b111111111111;
assign Lowerletter[4] = 12'b111111111111;
assign Lowerletter[5] = 12'b111111111111;
assign Lowerletter[6] = 12'b111111111111;
assign Lowerletter[7] = 12'b111111111111;
assign Lowerletter[8] = 12'b111111111111;
assign Lowerletter[9] = 12'b111111111111;
assign Lowerletter[10] = 12'b111111111111;
assign Lowerletter[11] = 12'b111111111111;
assign Lowerletter[12] = 12'b111111111111;
assign Lowerletter[13] = 12'b111111111111;
assign Lowerletter[14] = 12'b111111111111;
assign Lowerletter[15] = 12'b111111111111;
assign Lowerletter[16] = 12'b111111111111;
assign Lowerletter[17] = 12'b111111111111;
assign Lowerletter[18] = 12'b000000000000;
assign Lowerletter[19] = 12'b000000000000;
assign Lowerletter[20] = 12'b000000000000;
assign Lowerletter[21] = 12'b111111111111;
assign Lowerletter[22] = 12'b111111111111;
assign Lowerletter[23] = 12'b111111111111;
assign Lowerletter[24] = 12'b111111111111;
assign Lowerletter[25] = 12'b111111111111;
assign Lowerletter[26] = 12'b111111111111;
assign Lowerletter[27] = 12'b111111111111;
assign Lowerletter[28] = 12'b111111111111;
assign Lowerletter[29] = 12'b000000000000;
assign Lowerletter[30] = 12'b111111111111;
assign Lowerletter[31] = 12'b111111111111;
assign Lowerletter[32] = 12'b111111111111;
assign Lowerletter[33] = 12'b111111111111;
assign Lowerletter[34] = 12'b111111111111;
assign Lowerletter[35] = 12'b000000000000;
assign Lowerletter[36] = 12'b000000000000;
assign Lowerletter[37] = 12'b000000000000;
assign Lowerletter[38] = 12'b111111111111;
assign Lowerletter[39] = 12'b111111111111;
assign Lowerletter[40] = 12'b111111111111;
assign Lowerletter[41] = 12'b111111111111;
assign Lowerletter[42] = 12'b000000000000;
assign Lowerletter[43] = 12'b111111111111;
assign Lowerletter[44] = 12'b111111111111;
assign Lowerletter[45] = 12'b000000000000;
assign Lowerletter[46] = 12'b111111111111;
assign Lowerletter[47] = 12'b111111111111;
assign Lowerletter[48] = 12'b111111111111;
assign Lowerletter[49] = 12'b111111111111;
assign Lowerletter[50] = 12'b111111111111;
assign Lowerletter[51] = 12'b000000000000;
assign Lowerletter[52] = 12'b000000000000;
assign Lowerletter[53] = 12'b000000000000;
assign Lowerletter[54] = 12'b111111111111;
assign Lowerletter[55] = 12'b111111111111;
assign Lowerletter[56] = 12'b111111111111;
assign Lowerletter[57] = 12'b111111111111;
assign Lowerletter[58] = 12'b111111111111;
assign Lowerletter[59] = 12'b111111111111;
assign Lowerletter[60] = 12'b111111111111;
assign Lowerletter[61] = 12'b111111111111;
assign Lowerletter[62] = 12'b111111111111;
assign Lowerletter[63] = 12'b111111111111;
assign Lowerletter[64] = 12'b111111111111;
assign Lowerletter[65] = 12'b111111111111;
assign Lowerletter[66] = 12'b000000000000;
assign Lowerletter[67] = 12'b111111111111;
assign Lowerletter[68] = 12'b111111111111;
assign Lowerletter[69] = 12'b111111111111;
assign Lowerletter[70] = 12'b111111111111;
assign Lowerletter[71] = 12'b111111111111;
assign Lowerletter[72] = 12'b111111111111;
assign Lowerletter[73] = 12'b111111111111;
assign Lowerletter[74] = 12'b000000000000;
assign Lowerletter[75] = 12'b111111111111;
assign Lowerletter[76] = 12'b111111111111;
assign Lowerletter[77] = 12'b111111111111;
assign Lowerletter[78] = 12'b111111111111;
assign Lowerletter[79] = 12'b111111111111;
assign Lowerletter[80] = 12'b111111111111;
assign Lowerletter[81] = 12'b111111111111;
assign Lowerletter[82] = 12'b000000000000;
assign Lowerletter[83] = 12'b111111111111;
assign Lowerletter[84] = 12'b111111111111;
assign Lowerletter[85] = 12'b111111111111;
assign Lowerletter[86] = 12'b111111111111;
assign Lowerletter[87] = 12'b111111111111;
assign Lowerletter[88] = 12'b111111111111;
assign Lowerletter[89] = 12'b111111111111;
assign Lowerletter[90] = 12'b000000000000;
assign Lowerletter[91] = 12'b111111111111;
assign Lowerletter[92] = 12'b000000000000;
assign Lowerletter[93] = 12'b111111111111;
assign Lowerletter[94] = 12'b111111111111;
assign Lowerletter[95] = 12'b111111111111;
assign Lowerletter[96] = 12'b111111111111;
assign Lowerletter[97] = 12'b111111111111;
assign Lowerletter[98] = 12'b000000000000;
assign Lowerletter[99] = 12'b000000000000;
assign Lowerletter[100] = 12'b111111111111;
assign Lowerletter[101] = 12'b000000000000;
assign Lowerletter[102] = 12'b111111111111;
assign Lowerletter[103] = 12'b111111111111;
assign Lowerletter[104] = 12'b111111111111;
assign Lowerletter[105] = 12'b111111111111;
assign Lowerletter[106] = 12'b000000000000;
assign Lowerletter[107] = 12'b111111111111;
assign Lowerletter[108] = 12'b111111111111;
assign Lowerletter[109] = 12'b000000000000;
assign Lowerletter[110] = 12'b111111111111;
assign Lowerletter[111] = 12'b111111111111;
assign Lowerletter[112] = 12'b111111111111;
assign Lowerletter[113] = 12'b111111111111;
assign Lowerletter[114] = 12'b000000000000;
assign Lowerletter[115] = 12'b000000000000;
assign Lowerletter[116] = 12'b000000000000;
assign Lowerletter[117] = 12'b111111111111;
assign Lowerletter[118] = 12'b111111111111;
assign Lowerletter[119] = 12'b111111111111;
assign Lowerletter[120] = 12'b111111111111;
assign Lowerletter[121] = 12'b111111111111;
assign Lowerletter[122] = 12'b111111111111;
assign Lowerletter[123] = 12'b111111111111;
assign Lowerletter[124] = 12'b111111111111;
assign Lowerletter[125] = 12'b111111111111;
assign Lowerletter[126] = 12'b111111111111;
assign Lowerletter[127] = 12'b111111111111;
assign Lowerletter[128] = 12'b111111111111;
assign Lowerletter[129] = 12'b111111111111;
assign Lowerletter[130] = 12'b111111111111;
assign Lowerletter[131] = 12'b111111111111;
assign Lowerletter[132] = 12'b111111111111;
assign Lowerletter[133] = 12'b111111111111;
assign Lowerletter[134] = 12'b111111111111;
assign Lowerletter[135] = 12'b111111111111;
assign Lowerletter[136] = 12'b111111111111;
assign Lowerletter[137] = 12'b111111111111;
assign Lowerletter[138] = 12'b111111111111;
assign Lowerletter[139] = 12'b111111111111;
assign Lowerletter[140] = 12'b111111111111;
assign Lowerletter[141] = 12'b111111111111;
assign Lowerletter[142] = 12'b111111111111;
assign Lowerletter[143] = 12'b111111111111;
assign Lowerletter[144] = 12'b111111111111;
assign Lowerletter[145] = 12'b111111111111;
assign Lowerletter[146] = 12'b111111111111;
assign Lowerletter[147] = 12'b000000000000;
assign Lowerletter[148] = 12'b000000000000;
assign Lowerletter[149] = 12'b111111111111;
assign Lowerletter[150] = 12'b111111111111;
assign Lowerletter[151] = 12'b111111111111;
assign Lowerletter[152] = 12'b111111111111;
assign Lowerletter[153] = 12'b111111111111;
assign Lowerletter[154] = 12'b000000000000;
assign Lowerletter[155] = 12'b111111111111;
assign Lowerletter[156] = 12'b111111111111;
assign Lowerletter[157] = 12'b000000000000;
assign Lowerletter[158] = 12'b111111111111;
assign Lowerletter[159] = 12'b111111111111;
assign Lowerletter[160] = 12'b111111111111;
assign Lowerletter[161] = 12'b111111111111;
assign Lowerletter[162] = 12'b000000000000;
assign Lowerletter[163] = 12'b111111111111;
assign Lowerletter[164] = 12'b111111111111;
assign Lowerletter[165] = 12'b111111111111;
assign Lowerletter[166] = 12'b111111111111;
assign Lowerletter[167] = 12'b111111111111;
assign Lowerletter[168] = 12'b111111111111;
assign Lowerletter[169] = 12'b111111111111;
assign Lowerletter[170] = 12'b000000000000;
assign Lowerletter[171] = 12'b111111111111;
assign Lowerletter[172] = 12'b111111111111;
assign Lowerletter[173] = 12'b000000000000;
assign Lowerletter[174] = 12'b111111111111;
assign Lowerletter[175] = 12'b111111111111;
assign Lowerletter[176] = 12'b111111111111;
assign Lowerletter[177] = 12'b111111111111;
assign Lowerletter[178] = 12'b111111111111;
assign Lowerletter[179] = 12'b000000000000;
assign Lowerletter[180] = 12'b000000000000;
assign Lowerletter[181] = 12'b111111111111;
assign Lowerletter[182] = 12'b111111111111;
assign Lowerletter[183] = 12'b111111111111;
assign Lowerletter[184] = 12'b111111111111;
assign Lowerletter[185] = 12'b111111111111;
assign Lowerletter[186] = 12'b111111111111;
assign Lowerletter[187] = 12'b111111111111;
assign Lowerletter[188] = 12'b111111111111;
assign Lowerletter[189] = 12'b111111111111;
assign Lowerletter[190] = 12'b111111111111;
assign Lowerletter[191] = 12'b111111111111;
assign Lowerletter[192] = 12'b111111111111;
assign Lowerletter[193] = 12'b111111111111;
assign Lowerletter[194] = 12'b111111111111;
assign Lowerletter[195] = 12'b111111111111;
assign Lowerletter[196] = 12'b111111111111;
assign Lowerletter[197] = 12'b000000000000;
assign Lowerletter[198] = 12'b111111111111;
assign Lowerletter[199] = 12'b111111111111;
assign Lowerletter[200] = 12'b111111111111;
assign Lowerletter[201] = 12'b111111111111;
assign Lowerletter[202] = 12'b111111111111;
assign Lowerletter[203] = 12'b111111111111;
assign Lowerletter[204] = 12'b111111111111;
assign Lowerletter[205] = 12'b000000000000;
assign Lowerletter[206] = 12'b111111111111;
assign Lowerletter[207] = 12'b111111111111;
assign Lowerletter[208] = 12'b111111111111;
assign Lowerletter[209] = 12'b111111111111;
assign Lowerletter[210] = 12'b111111111111;
assign Lowerletter[211] = 12'b111111111111;
assign Lowerletter[212] = 12'b111111111111;
assign Lowerletter[213] = 12'b000000000000;
assign Lowerletter[214] = 12'b111111111111;
assign Lowerletter[215] = 12'b111111111111;
assign Lowerletter[216] = 12'b111111111111;
assign Lowerletter[217] = 12'b111111111111;
assign Lowerletter[218] = 12'b111111111111;
assign Lowerletter[219] = 12'b000000000000;
assign Lowerletter[220] = 12'b000000000000;
assign Lowerletter[221] = 12'b000000000000;
assign Lowerletter[222] = 12'b111111111111;
assign Lowerletter[223] = 12'b111111111111;
assign Lowerletter[224] = 12'b111111111111;
assign Lowerletter[225] = 12'b111111111111;
assign Lowerletter[226] = 12'b000000000000;
assign Lowerletter[227] = 12'b111111111111;
assign Lowerletter[228] = 12'b111111111111;
assign Lowerletter[229] = 12'b000000000000;
assign Lowerletter[230] = 12'b111111111111;
assign Lowerletter[231] = 12'b111111111111;
assign Lowerletter[232] = 12'b111111111111;
assign Lowerletter[233] = 12'b111111111111;
assign Lowerletter[234] = 12'b000000000000;
assign Lowerletter[235] = 12'b111111111111;
assign Lowerletter[236] = 12'b111111111111;
assign Lowerletter[237] = 12'b000000000000;
assign Lowerletter[238] = 12'b111111111111;
assign Lowerletter[239] = 12'b111111111111;
assign Lowerletter[240] = 12'b111111111111;
assign Lowerletter[241] = 12'b111111111111;
assign Lowerletter[242] = 12'b000000000000;
assign Lowerletter[243] = 12'b000000000000;
assign Lowerletter[244] = 12'b000000000000;
assign Lowerletter[245] = 12'b000000000000;
assign Lowerletter[246] = 12'b111111111111;
assign Lowerletter[247] = 12'b111111111111;
assign Lowerletter[248] = 12'b111111111111;
assign Lowerletter[249] = 12'b111111111111;
assign Lowerletter[250] = 12'b111111111111;
assign Lowerletter[251] = 12'b111111111111;
assign Lowerletter[252] = 12'b111111111111;
assign Lowerletter[253] = 12'b111111111111;
assign Lowerletter[254] = 12'b111111111111;
assign Lowerletter[255] = 12'b111111111111;
assign Lowerletter[256] = 12'b111111111111;
assign Lowerletter[257] = 12'b111111111111;
assign Lowerletter[258] = 12'b111111111111;
assign Lowerletter[259] = 12'b111111111111;
assign Lowerletter[260] = 12'b111111111111;
assign Lowerletter[261] = 12'b111111111111;
assign Lowerletter[262] = 12'b111111111111;
assign Lowerletter[263] = 12'b111111111111;
assign Lowerletter[264] = 12'b111111111111;
assign Lowerletter[265] = 12'b111111111111;
assign Lowerletter[266] = 12'b111111111111;
assign Lowerletter[267] = 12'b111111111111;
assign Lowerletter[268] = 12'b111111111111;
assign Lowerletter[269] = 12'b111111111111;
assign Lowerletter[270] = 12'b111111111111;
assign Lowerletter[271] = 12'b111111111111;
assign Lowerletter[272] = 12'b111111111111;
assign Lowerletter[273] = 12'b111111111111;
assign Lowerletter[274] = 12'b111111111111;
assign Lowerletter[275] = 12'b000000000000;
assign Lowerletter[276] = 12'b000000000000;
assign Lowerletter[277] = 12'b000000000000;
assign Lowerletter[278] = 12'b111111111111;
assign Lowerletter[279] = 12'b111111111111;
assign Lowerletter[280] = 12'b111111111111;
assign Lowerletter[281] = 12'b111111111111;
assign Lowerletter[282] = 12'b000000000000;
assign Lowerletter[283] = 12'b111111111111;
assign Lowerletter[284] = 12'b111111111111;
assign Lowerletter[285] = 12'b000000000000;
assign Lowerletter[286] = 12'b111111111111;
assign Lowerletter[287] = 12'b111111111111;
assign Lowerletter[288] = 12'b111111111111;
assign Lowerletter[289] = 12'b111111111111;
assign Lowerletter[290] = 12'b000000000000;
assign Lowerletter[291] = 12'b000000000000;
assign Lowerletter[292] = 12'b000000000000;
assign Lowerletter[293] = 12'b111111111111;
assign Lowerletter[294] = 12'b111111111111;
assign Lowerletter[295] = 12'b111111111111;
assign Lowerletter[296] = 12'b111111111111;
assign Lowerletter[297] = 12'b111111111111;
assign Lowerletter[298] = 12'b000000000000;
assign Lowerletter[299] = 12'b111111111111;
assign Lowerletter[300] = 12'b111111111111;
assign Lowerletter[301] = 12'b111111111111;
assign Lowerletter[302] = 12'b111111111111;
assign Lowerletter[303] = 12'b111111111111;
assign Lowerletter[304] = 12'b111111111111;
assign Lowerletter[305] = 12'b111111111111;
assign Lowerletter[306] = 12'b111111111111;
assign Lowerletter[307] = 12'b000000000000;
assign Lowerletter[308] = 12'b000000000000;
assign Lowerletter[309] = 12'b000000000000;
assign Lowerletter[310] = 12'b111111111111;
assign Lowerletter[311] = 12'b111111111111;
assign Lowerletter[312] = 12'b111111111111;
assign Lowerletter[313] = 12'b111111111111;
assign Lowerletter[314] = 12'b111111111111;
assign Lowerletter[315] = 12'b111111111111;
assign Lowerletter[316] = 12'b111111111111;
assign Lowerletter[317] = 12'b111111111111;
assign Lowerletter[318] = 12'b111111111111;
assign Lowerletter[319] = 12'b111111111111;
assign Lowerletter[320] = 12'b111111111111;
assign Lowerletter[321] = 12'b111111111111;
assign Lowerletter[322] = 12'b111111111111;
assign Lowerletter[323] = 12'b000000000000;
assign Lowerletter[324] = 12'b000000000000;
assign Lowerletter[325] = 12'b111111111111;
assign Lowerletter[326] = 12'b111111111111;
assign Lowerletter[327] = 12'b111111111111;
assign Lowerletter[328] = 12'b111111111111;
assign Lowerletter[329] = 12'b111111111111;
assign Lowerletter[330] = 12'b111111111111;
assign Lowerletter[331] = 12'b000000000000;
assign Lowerletter[332] = 12'b111111111111;
assign Lowerletter[333] = 12'b111111111111;
assign Lowerletter[334] = 12'b111111111111;
assign Lowerletter[335] = 12'b111111111111;
assign Lowerletter[336] = 12'b111111111111;
assign Lowerletter[337] = 12'b111111111111;
assign Lowerletter[338] = 12'b000000000000;
assign Lowerletter[339] = 12'b000000000000;
assign Lowerletter[340] = 12'b000000000000;
assign Lowerletter[341] = 12'b000000000000;
assign Lowerletter[342] = 12'b111111111111;
assign Lowerletter[343] = 12'b111111111111;
assign Lowerletter[344] = 12'b111111111111;
assign Lowerletter[345] = 12'b111111111111;
assign Lowerletter[346] = 12'b111111111111;
assign Lowerletter[347] = 12'b000000000000;
assign Lowerletter[348] = 12'b111111111111;
assign Lowerletter[349] = 12'b111111111111;
assign Lowerletter[350] = 12'b111111111111;
assign Lowerletter[351] = 12'b111111111111;
assign Lowerletter[352] = 12'b111111111111;
assign Lowerletter[353] = 12'b111111111111;
assign Lowerletter[354] = 12'b111111111111;
assign Lowerletter[355] = 12'b000000000000;
assign Lowerletter[356] = 12'b111111111111;
assign Lowerletter[357] = 12'b111111111111;
assign Lowerletter[358] = 12'b111111111111;
assign Lowerletter[359] = 12'b111111111111;
assign Lowerletter[360] = 12'b111111111111;
assign Lowerletter[361] = 12'b111111111111;
assign Lowerletter[362] = 12'b111111111111;
assign Lowerletter[363] = 12'b000000000000;
assign Lowerletter[364] = 12'b111111111111;
assign Lowerletter[365] = 12'b111111111111;
assign Lowerletter[366] = 12'b111111111111;
assign Lowerletter[367] = 12'b111111111111;
assign Lowerletter[368] = 12'b111111111111;
assign Lowerletter[369] = 12'b111111111111;
assign Lowerletter[370] = 12'b111111111111;
assign Lowerletter[371] = 12'b000000000000;
assign Lowerletter[372] = 12'b111111111111;
assign Lowerletter[373] = 12'b111111111111;
assign Lowerletter[374] = 12'b111111111111;
assign Lowerletter[375] = 12'b111111111111;
assign Lowerletter[376] = 12'b111111111111;
assign Lowerletter[377] = 12'b111111111111;
assign Lowerletter[378] = 12'b111111111111;
assign Lowerletter[379] = 12'b111111111111;
assign Lowerletter[380] = 12'b111111111111;
assign Lowerletter[381] = 12'b111111111111;
assign Lowerletter[382] = 12'b111111111111;
assign Lowerletter[383] = 12'b111111111111;
assign Lowerletter[384] = 12'b111111111111;
assign Lowerletter[385] = 12'b111111111111;
assign Lowerletter[386] = 12'b111111111111;
assign Lowerletter[387] = 12'b111111111111;
assign Lowerletter[388] = 12'b111111111111;
assign Lowerletter[389] = 12'b111111111111;
assign Lowerletter[390] = 12'b111111111111;
assign Lowerletter[391] = 12'b111111111111;
assign Lowerletter[392] = 12'b111111111111;
assign Lowerletter[393] = 12'b111111111111;
assign Lowerletter[394] = 12'b111111111111;
assign Lowerletter[395] = 12'b111111111111;
assign Lowerletter[396] = 12'b111111111111;
assign Lowerletter[397] = 12'b111111111111;
assign Lowerletter[398] = 12'b111111111111;
assign Lowerletter[399] = 12'b111111111111;
assign Lowerletter[400] = 12'b111111111111;
assign Lowerletter[401] = 12'b111111111111;
assign Lowerletter[402] = 12'b111111111111;
assign Lowerletter[403] = 12'b000000000000;
assign Lowerletter[404] = 12'b000000000000;
assign Lowerletter[405] = 12'b000000000000;
assign Lowerletter[406] = 12'b111111111111;
assign Lowerletter[407] = 12'b111111111111;
assign Lowerletter[408] = 12'b111111111111;
assign Lowerletter[409] = 12'b111111111111;
assign Lowerletter[410] = 12'b000000000000;
assign Lowerletter[411] = 12'b111111111111;
assign Lowerletter[412] = 12'b111111111111;
assign Lowerletter[413] = 12'b000000000000;
assign Lowerletter[414] = 12'b111111111111;
assign Lowerletter[415] = 12'b111111111111;
assign Lowerletter[416] = 12'b111111111111;
assign Lowerletter[417] = 12'b111111111111;
assign Lowerletter[418] = 12'b111111111111;
assign Lowerletter[419] = 12'b000000000000;
assign Lowerletter[420] = 12'b000000000000;
assign Lowerletter[421] = 12'b000000000000;
assign Lowerletter[422] = 12'b111111111111;
assign Lowerletter[423] = 12'b111111111111;
assign Lowerletter[424] = 12'b111111111111;
assign Lowerletter[425] = 12'b111111111111;
assign Lowerletter[426] = 12'b111111111111;
assign Lowerletter[427] = 12'b111111111111;
assign Lowerletter[428] = 12'b111111111111;
assign Lowerletter[429] = 12'b000000000000;
assign Lowerletter[430] = 12'b111111111111;
assign Lowerletter[431] = 12'b111111111111;
assign Lowerletter[432] = 12'b111111111111;
assign Lowerletter[433] = 12'b111111111111;
assign Lowerletter[434] = 12'b000000000000;
assign Lowerletter[435] = 12'b111111111111;
assign Lowerletter[436] = 12'b111111111111;
assign Lowerletter[437] = 12'b000000000000;
assign Lowerletter[438] = 12'b111111111111;
assign Lowerletter[439] = 12'b111111111111;
assign Lowerletter[440] = 12'b111111111111;
assign Lowerletter[441] = 12'b111111111111;
assign Lowerletter[442] = 12'b111111111111;
assign Lowerletter[443] = 12'b000000000000;
assign Lowerletter[444] = 12'b000000000000;
assign Lowerletter[445] = 12'b111111111111;
assign Lowerletter[446] = 12'b111111111111;
assign Lowerletter[447] = 12'b111111111111;
assign Lowerletter[448] = 12'b111111111111;
assign Lowerletter[449] = 12'b111111111111;
assign Lowerletter[450] = 12'b000000000000;
assign Lowerletter[451] = 12'b111111111111;
assign Lowerletter[452] = 12'b111111111111;
assign Lowerletter[453] = 12'b111111111111;
assign Lowerletter[454] = 12'b111111111111;
assign Lowerletter[455] = 12'b111111111111;
assign Lowerletter[456] = 12'b111111111111;
assign Lowerletter[457] = 12'b111111111111;
assign Lowerletter[458] = 12'b000000000000;
assign Lowerletter[459] = 12'b111111111111;
assign Lowerletter[460] = 12'b111111111111;
assign Lowerletter[461] = 12'b111111111111;
assign Lowerletter[462] = 12'b111111111111;
assign Lowerletter[463] = 12'b111111111111;
assign Lowerletter[464] = 12'b111111111111;
assign Lowerletter[465] = 12'b111111111111;
assign Lowerletter[466] = 12'b000000000000;
assign Lowerletter[467] = 12'b111111111111;
assign Lowerletter[468] = 12'b111111111111;
assign Lowerletter[469] = 12'b111111111111;
assign Lowerletter[470] = 12'b111111111111;
assign Lowerletter[471] = 12'b111111111111;
assign Lowerletter[472] = 12'b111111111111;
assign Lowerletter[473] = 12'b111111111111;
assign Lowerletter[474] = 12'b000000000000;
assign Lowerletter[475] = 12'b111111111111;
assign Lowerletter[476] = 12'b000000000000;
assign Lowerletter[477] = 12'b111111111111;
assign Lowerletter[478] = 12'b111111111111;
assign Lowerletter[479] = 12'b111111111111;
assign Lowerletter[480] = 12'b111111111111;
assign Lowerletter[481] = 12'b111111111111;
assign Lowerletter[482] = 12'b000000000000;
assign Lowerletter[483] = 12'b000000000000;
assign Lowerletter[484] = 12'b111111111111;
assign Lowerletter[485] = 12'b000000000000;
assign Lowerletter[486] = 12'b111111111111;
assign Lowerletter[487] = 12'b111111111111;
assign Lowerletter[488] = 12'b111111111111;
assign Lowerletter[489] = 12'b111111111111;
assign Lowerletter[490] = 12'b000000000000;
assign Lowerletter[491] = 12'b111111111111;
assign Lowerletter[492] = 12'b111111111111;
assign Lowerletter[493] = 12'b000000000000;
assign Lowerletter[494] = 12'b111111111111;
assign Lowerletter[495] = 12'b111111111111;
assign Lowerletter[496] = 12'b111111111111;
assign Lowerletter[497] = 12'b111111111111;
assign Lowerletter[498] = 12'b000000000000;
assign Lowerletter[499] = 12'b111111111111;
assign Lowerletter[500] = 12'b111111111111;
assign Lowerletter[501] = 12'b000000000000;
assign Lowerletter[502] = 12'b111111111111;
assign Lowerletter[503] = 12'b111111111111;
assign Lowerletter[504] = 12'b111111111111;
assign Lowerletter[505] = 12'b111111111111;
assign Lowerletter[506] = 12'b111111111111;
assign Lowerletter[507] = 12'b111111111111;
assign Lowerletter[508] = 12'b111111111111;
assign Lowerletter[509] = 12'b111111111111;
assign Lowerletter[510] = 12'b111111111111;
assign Lowerletter[511] = 12'b111111111111;
assign Lowerletter[512] = 12'b111111111111;
assign Lowerletter[513] = 12'b111111111111;
assign Lowerletter[514] = 12'b111111111111;
assign Lowerletter[515] = 12'b111111111111;
assign Lowerletter[516] = 12'b111111111111;
assign Lowerletter[517] = 12'b111111111111;
assign Lowerletter[518] = 12'b111111111111;
assign Lowerletter[519] = 12'b111111111111;
assign Lowerletter[520] = 12'b111111111111;
assign Lowerletter[521] = 12'b111111111111;
assign Lowerletter[522] = 12'b111111111111;
assign Lowerletter[523] = 12'b000000000000;
assign Lowerletter[524] = 12'b111111111111;
assign Lowerletter[525] = 12'b111111111111;
assign Lowerletter[526] = 12'b111111111111;
assign Lowerletter[527] = 12'b111111111111;
assign Lowerletter[528] = 12'b111111111111;
assign Lowerletter[529] = 12'b111111111111;
assign Lowerletter[530] = 12'b111111111111;
assign Lowerletter[531] = 12'b111111111111;
assign Lowerletter[532] = 12'b111111111111;
assign Lowerletter[533] = 12'b111111111111;
assign Lowerletter[534] = 12'b111111111111;
assign Lowerletter[535] = 12'b111111111111;
assign Lowerletter[536] = 12'b111111111111;
assign Lowerletter[537] = 12'b111111111111;
assign Lowerletter[538] = 12'b111111111111;
assign Lowerletter[539] = 12'b000000000000;
assign Lowerletter[540] = 12'b111111111111;
assign Lowerletter[541] = 12'b111111111111;
assign Lowerletter[542] = 12'b111111111111;
assign Lowerletter[543] = 12'b111111111111;
assign Lowerletter[544] = 12'b111111111111;
assign Lowerletter[545] = 12'b111111111111;
assign Lowerletter[546] = 12'b111111111111;
assign Lowerletter[547] = 12'b000000000000;
assign Lowerletter[548] = 12'b111111111111;
assign Lowerletter[549] = 12'b111111111111;
assign Lowerletter[550] = 12'b111111111111;
assign Lowerletter[551] = 12'b111111111111;
assign Lowerletter[552] = 12'b111111111111;
assign Lowerletter[553] = 12'b111111111111;
assign Lowerletter[554] = 12'b111111111111;
assign Lowerletter[555] = 12'b000000000000;
assign Lowerletter[556] = 12'b111111111111;
assign Lowerletter[557] = 12'b111111111111;
assign Lowerletter[558] = 12'b111111111111;
assign Lowerletter[559] = 12'b111111111111;
assign Lowerletter[560] = 12'b111111111111;
assign Lowerletter[561] = 12'b111111111111;
assign Lowerletter[562] = 12'b111111111111;
assign Lowerletter[563] = 12'b000000000000;
assign Lowerletter[564] = 12'b111111111111;
assign Lowerletter[565] = 12'b111111111111;
assign Lowerletter[566] = 12'b111111111111;
assign Lowerletter[567] = 12'b111111111111;
assign Lowerletter[568] = 12'b111111111111;
assign Lowerletter[569] = 12'b111111111111;
assign Lowerletter[570] = 12'b111111111111;
assign Lowerletter[571] = 12'b111111111111;
assign Lowerletter[572] = 12'b111111111111;
assign Lowerletter[573] = 12'b111111111111;
assign Lowerletter[574] = 12'b111111111111;
assign Lowerletter[575] = 12'b111111111111;
assign Lowerletter[576] = 12'b111111111111;
assign Lowerletter[577] = 12'b111111111111;
assign Lowerletter[578] = 12'b111111111111;
assign Lowerletter[579] = 12'b111111111111;
assign Lowerletter[580] = 12'b111111111111;
assign Lowerletter[581] = 12'b111111111111;
assign Lowerletter[582] = 12'b111111111111;
assign Lowerletter[583] = 12'b111111111111;
assign Lowerletter[584] = 12'b111111111111;
assign Lowerletter[585] = 12'b111111111111;
assign Lowerletter[586] = 12'b111111111111;
assign Lowerletter[587] = 12'b111111111111;
assign Lowerletter[588] = 12'b111111111111;
assign Lowerletter[589] = 12'b111111111111;
assign Lowerletter[590] = 12'b111111111111;
assign Lowerletter[591] = 12'b111111111111;
assign Lowerletter[592] = 12'b111111111111;
assign Lowerletter[593] = 12'b111111111111;
assign Lowerletter[594] = 12'b111111111111;
assign Lowerletter[595] = 12'b111111111111;
assign Lowerletter[596] = 12'b000000000000;
assign Lowerletter[597] = 12'b111111111111;
assign Lowerletter[598] = 12'b111111111111;
assign Lowerletter[599] = 12'b111111111111;
assign Lowerletter[600] = 12'b111111111111;
assign Lowerletter[601] = 12'b111111111111;
assign Lowerletter[602] = 12'b111111111111;
assign Lowerletter[603] = 12'b111111111111;
assign Lowerletter[604] = 12'b111111111111;
assign Lowerletter[605] = 12'b111111111111;
assign Lowerletter[606] = 12'b111111111111;
assign Lowerletter[607] = 12'b111111111111;
assign Lowerletter[608] = 12'b111111111111;
assign Lowerletter[609] = 12'b111111111111;
assign Lowerletter[610] = 12'b111111111111;
assign Lowerletter[611] = 12'b111111111111;
assign Lowerletter[612] = 12'b000000000000;
assign Lowerletter[613] = 12'b111111111111;
assign Lowerletter[614] = 12'b111111111111;
assign Lowerletter[615] = 12'b111111111111;
assign Lowerletter[616] = 12'b111111111111;
assign Lowerletter[617] = 12'b111111111111;
assign Lowerletter[618] = 12'b111111111111;
assign Lowerletter[619] = 12'b111111111111;
assign Lowerletter[620] = 12'b000000000000;
assign Lowerletter[621] = 12'b111111111111;
assign Lowerletter[622] = 12'b111111111111;
assign Lowerletter[623] = 12'b111111111111;
assign Lowerletter[624] = 12'b111111111111;
assign Lowerletter[625] = 12'b111111111111;
assign Lowerletter[626] = 12'b000000000000;
assign Lowerletter[627] = 12'b111111111111;
assign Lowerletter[628] = 12'b000000000000;
assign Lowerletter[629] = 12'b111111111111;
assign Lowerletter[630] = 12'b111111111111;
assign Lowerletter[631] = 12'b111111111111;
assign Lowerletter[632] = 12'b111111111111;
assign Lowerletter[633] = 12'b111111111111;
assign Lowerletter[634] = 12'b111111111111;
assign Lowerletter[635] = 12'b000000000000;
assign Lowerletter[636] = 12'b111111111111;
assign Lowerletter[637] = 12'b111111111111;
assign Lowerletter[638] = 12'b111111111111;
assign Lowerletter[639] = 12'b111111111111;
assign Lowerletter[640] = 12'b111111111111;
assign Lowerletter[641] = 12'b111111111111;
assign Lowerletter[642] = 12'b000000000000;
assign Lowerletter[643] = 12'b111111111111;
assign Lowerletter[644] = 12'b111111111111;
assign Lowerletter[645] = 12'b111111111111;
assign Lowerletter[646] = 12'b111111111111;
assign Lowerletter[647] = 12'b111111111111;
assign Lowerletter[648] = 12'b111111111111;
assign Lowerletter[649] = 12'b111111111111;
assign Lowerletter[650] = 12'b000000000000;
assign Lowerletter[651] = 12'b111111111111;
assign Lowerletter[652] = 12'b111111111111;
assign Lowerletter[653] = 12'b111111111111;
assign Lowerletter[654] = 12'b111111111111;
assign Lowerletter[655] = 12'b111111111111;
assign Lowerletter[656] = 12'b111111111111;
assign Lowerletter[657] = 12'b111111111111;
assign Lowerletter[658] = 12'b000000000000;
assign Lowerletter[659] = 12'b111111111111;
assign Lowerletter[660] = 12'b111111111111;
assign Lowerletter[661] = 12'b000000000000;
assign Lowerletter[662] = 12'b111111111111;
assign Lowerletter[663] = 12'b111111111111;
assign Lowerletter[664] = 12'b111111111111;
assign Lowerletter[665] = 12'b111111111111;
assign Lowerletter[666] = 12'b000000000000;
assign Lowerletter[667] = 12'b111111111111;
assign Lowerletter[668] = 12'b000000000000;
assign Lowerletter[669] = 12'b111111111111;
assign Lowerletter[670] = 12'b111111111111;
assign Lowerletter[671] = 12'b111111111111;
assign Lowerletter[672] = 12'b111111111111;
assign Lowerletter[673] = 12'b111111111111;
assign Lowerletter[674] = 12'b000000000000;
assign Lowerletter[675] = 12'b000000000000;
assign Lowerletter[676] = 12'b111111111111;
assign Lowerletter[677] = 12'b111111111111;
assign Lowerletter[678] = 12'b111111111111;
assign Lowerletter[679] = 12'b111111111111;
assign Lowerletter[680] = 12'b111111111111;
assign Lowerletter[681] = 12'b111111111111;
assign Lowerletter[682] = 12'b000000000000;
assign Lowerletter[683] = 12'b111111111111;
assign Lowerletter[684] = 12'b000000000000;
assign Lowerletter[685] = 12'b111111111111;
assign Lowerletter[686] = 12'b111111111111;
assign Lowerletter[687] = 12'b111111111111;
assign Lowerletter[688] = 12'b111111111111;
assign Lowerletter[689] = 12'b111111111111;
assign Lowerletter[690] = 12'b000000000000;
assign Lowerletter[691] = 12'b111111111111;
assign Lowerletter[692] = 12'b111111111111;
assign Lowerletter[693] = 12'b000000000000;
assign Lowerletter[694] = 12'b111111111111;
assign Lowerletter[695] = 12'b111111111111;
assign Lowerletter[696] = 12'b111111111111;
assign Lowerletter[697] = 12'b111111111111;
assign Lowerletter[698] = 12'b111111111111;
assign Lowerletter[699] = 12'b111111111111;
assign Lowerletter[700] = 12'b111111111111;
assign Lowerletter[701] = 12'b111111111111;
assign Lowerletter[702] = 12'b111111111111;
assign Lowerletter[703] = 12'b111111111111;
assign Lowerletter[704] = 12'b111111111111;
assign Lowerletter[705] = 12'b111111111111;
assign Lowerletter[706] = 12'b111111111111;
assign Lowerletter[707] = 12'b000000000000;
assign Lowerletter[708] = 12'b111111111111;
assign Lowerletter[709] = 12'b111111111111;
assign Lowerletter[710] = 12'b111111111111;
assign Lowerletter[711] = 12'b111111111111;
assign Lowerletter[712] = 12'b111111111111;
assign Lowerletter[713] = 12'b111111111111;
assign Lowerletter[714] = 12'b111111111111;
assign Lowerletter[715] = 12'b000000000000;
assign Lowerletter[716] = 12'b111111111111;
assign Lowerletter[717] = 12'b111111111111;
assign Lowerletter[718] = 12'b111111111111;
assign Lowerletter[719] = 12'b111111111111;
assign Lowerletter[720] = 12'b111111111111;
assign Lowerletter[721] = 12'b111111111111;
assign Lowerletter[722] = 12'b111111111111;
assign Lowerletter[723] = 12'b000000000000;
assign Lowerletter[724] = 12'b111111111111;
assign Lowerletter[725] = 12'b111111111111;
assign Lowerletter[726] = 12'b111111111111;
assign Lowerletter[727] = 12'b111111111111;
assign Lowerletter[728] = 12'b111111111111;
assign Lowerletter[729] = 12'b111111111111;
assign Lowerletter[730] = 12'b111111111111;
assign Lowerletter[731] = 12'b000000000000;
assign Lowerletter[732] = 12'b111111111111;
assign Lowerletter[733] = 12'b111111111111;
assign Lowerletter[734] = 12'b111111111111;
assign Lowerletter[735] = 12'b111111111111;
assign Lowerletter[736] = 12'b111111111111;
assign Lowerletter[737] = 12'b111111111111;
assign Lowerletter[738] = 12'b111111111111;
assign Lowerletter[739] = 12'b000000000000;
assign Lowerletter[740] = 12'b111111111111;
assign Lowerletter[741] = 12'b111111111111;
assign Lowerletter[742] = 12'b111111111111;
assign Lowerletter[743] = 12'b111111111111;
assign Lowerletter[744] = 12'b111111111111;
assign Lowerletter[745] = 12'b111111111111;
assign Lowerletter[746] = 12'b111111111111;
assign Lowerletter[747] = 12'b000000000000;
assign Lowerletter[748] = 12'b111111111111;
assign Lowerletter[749] = 12'b111111111111;
assign Lowerletter[750] = 12'b111111111111;
assign Lowerletter[751] = 12'b111111111111;
assign Lowerletter[752] = 12'b111111111111;
assign Lowerletter[753] = 12'b111111111111;
assign Lowerletter[754] = 12'b111111111111;
assign Lowerletter[755] = 12'b000000000000;
assign Lowerletter[756] = 12'b111111111111;
assign Lowerletter[757] = 12'b111111111111;
assign Lowerletter[758] = 12'b111111111111;
assign Lowerletter[759] = 12'b111111111111;
assign Lowerletter[760] = 12'b111111111111;
assign Lowerletter[761] = 12'b111111111111;
assign Lowerletter[762] = 12'b111111111111;
assign Lowerletter[763] = 12'b111111111111;
assign Lowerletter[764] = 12'b111111111111;
assign Lowerletter[765] = 12'b111111111111;
assign Lowerletter[766] = 12'b111111111111;
assign Lowerletter[767] = 12'b111111111111;
assign Lowerletter[768] = 12'b111111111111;
assign Lowerletter[769] = 12'b111111111111;
assign Lowerletter[770] = 12'b111111111111;
assign Lowerletter[771] = 12'b111111111111;
assign Lowerletter[772] = 12'b111111111111;
assign Lowerletter[773] = 12'b111111111111;
assign Lowerletter[774] = 12'b111111111111;
assign Lowerletter[775] = 12'b111111111111;
assign Lowerletter[776] = 12'b111111111111;
assign Lowerletter[777] = 12'b111111111111;
assign Lowerletter[778] = 12'b111111111111;
assign Lowerletter[779] = 12'b111111111111;
assign Lowerletter[780] = 12'b111111111111;
assign Lowerletter[781] = 12'b111111111111;
assign Lowerletter[782] = 12'b111111111111;
assign Lowerletter[783] = 12'b111111111111;
assign Lowerletter[784] = 12'b111111111111;
assign Lowerletter[785] = 12'b000000000000;
assign Lowerletter[786] = 12'b000000000000;
assign Lowerletter[787] = 12'b111111111111;
assign Lowerletter[788] = 12'b000000000000;
assign Lowerletter[789] = 12'b111111111111;
assign Lowerletter[790] = 12'b111111111111;
assign Lowerletter[791] = 12'b111111111111;
assign Lowerletter[792] = 12'b111111111111;
assign Lowerletter[793] = 12'b000000000000;
assign Lowerletter[794] = 12'b111111111111;
assign Lowerletter[795] = 12'b000000000000;
assign Lowerletter[796] = 12'b111111111111;
assign Lowerletter[797] = 12'b000000000000;
assign Lowerletter[798] = 12'b111111111111;
assign Lowerletter[799] = 12'b111111111111;
assign Lowerletter[800] = 12'b111111111111;
assign Lowerletter[801] = 12'b000000000000;
assign Lowerletter[802] = 12'b111111111111;
assign Lowerletter[803] = 12'b000000000000;
assign Lowerletter[804] = 12'b111111111111;
assign Lowerletter[805] = 12'b000000000000;
assign Lowerletter[806] = 12'b111111111111;
assign Lowerletter[807] = 12'b111111111111;
assign Lowerletter[808] = 12'b111111111111;
assign Lowerletter[809] = 12'b000000000000;
assign Lowerletter[810] = 12'b111111111111;
assign Lowerletter[811] = 12'b000000000000;
assign Lowerletter[812] = 12'b111111111111;
assign Lowerletter[813] = 12'b000000000000;
assign Lowerletter[814] = 12'b111111111111;
assign Lowerletter[815] = 12'b111111111111;
assign Lowerletter[816] = 12'b111111111111;
assign Lowerletter[817] = 12'b000000000000;
assign Lowerletter[818] = 12'b111111111111;
assign Lowerletter[819] = 12'b000000000000;
assign Lowerletter[820] = 12'b111111111111;
assign Lowerletter[821] = 12'b000000000000;
assign Lowerletter[822] = 12'b111111111111;
assign Lowerletter[823] = 12'b111111111111;
assign Lowerletter[824] = 12'b111111111111;
assign Lowerletter[825] = 12'b111111111111;
assign Lowerletter[826] = 12'b111111111111;
assign Lowerletter[827] = 12'b111111111111;
assign Lowerletter[828] = 12'b111111111111;
assign Lowerletter[829] = 12'b111111111111;
assign Lowerletter[830] = 12'b111111111111;
assign Lowerletter[831] = 12'b111111111111;
assign Lowerletter[832] = 12'b111111111111;
assign Lowerletter[833] = 12'b111111111111;
assign Lowerletter[834] = 12'b111111111111;
assign Lowerletter[835] = 12'b111111111111;
assign Lowerletter[836] = 12'b111111111111;
assign Lowerletter[837] = 12'b111111111111;
assign Lowerletter[838] = 12'b111111111111;
assign Lowerletter[839] = 12'b111111111111;
assign Lowerletter[840] = 12'b111111111111;
assign Lowerletter[841] = 12'b111111111111;
assign Lowerletter[842] = 12'b111111111111;
assign Lowerletter[843] = 12'b111111111111;
assign Lowerletter[844] = 12'b111111111111;
assign Lowerletter[845] = 12'b111111111111;
assign Lowerletter[846] = 12'b111111111111;
assign Lowerletter[847] = 12'b111111111111;
assign Lowerletter[848] = 12'b111111111111;
assign Lowerletter[849] = 12'b111111111111;
assign Lowerletter[850] = 12'b000000000000;
assign Lowerletter[851] = 12'b000000000000;
assign Lowerletter[852] = 12'b000000000000;
assign Lowerletter[853] = 12'b111111111111;
assign Lowerletter[854] = 12'b111111111111;
assign Lowerletter[855] = 12'b111111111111;
assign Lowerletter[856] = 12'b111111111111;
assign Lowerletter[857] = 12'b111111111111;
assign Lowerletter[858] = 12'b000000000000;
assign Lowerletter[859] = 12'b111111111111;
assign Lowerletter[860] = 12'b111111111111;
assign Lowerletter[861] = 12'b000000000000;
assign Lowerletter[862] = 12'b111111111111;
assign Lowerletter[863] = 12'b111111111111;
assign Lowerletter[864] = 12'b111111111111;
assign Lowerletter[865] = 12'b111111111111;
assign Lowerletter[866] = 12'b000000000000;
assign Lowerletter[867] = 12'b111111111111;
assign Lowerletter[868] = 12'b111111111111;
assign Lowerletter[869] = 12'b000000000000;
assign Lowerletter[870] = 12'b111111111111;
assign Lowerletter[871] = 12'b111111111111;
assign Lowerletter[872] = 12'b111111111111;
assign Lowerletter[873] = 12'b111111111111;
assign Lowerletter[874] = 12'b000000000000;
assign Lowerletter[875] = 12'b111111111111;
assign Lowerletter[876] = 12'b111111111111;
assign Lowerletter[877] = 12'b000000000000;
assign Lowerletter[878] = 12'b111111111111;
assign Lowerletter[879] = 12'b111111111111;
assign Lowerletter[880] = 12'b111111111111;
assign Lowerletter[881] = 12'b111111111111;
assign Lowerletter[882] = 12'b000000000000;
assign Lowerletter[883] = 12'b111111111111;
assign Lowerletter[884] = 12'b111111111111;
assign Lowerletter[885] = 12'b000000000000;
assign Lowerletter[886] = 12'b111111111111;
assign Lowerletter[887] = 12'b111111111111;
assign Lowerletter[888] = 12'b111111111111;
assign Lowerletter[889] = 12'b111111111111;
assign Lowerletter[890] = 12'b111111111111;
assign Lowerletter[891] = 12'b111111111111;
assign Lowerletter[892] = 12'b111111111111;
assign Lowerletter[893] = 12'b111111111111;
assign Lowerletter[894] = 12'b111111111111;
assign Lowerletter[895] = 12'b111111111111;
assign Lowerletter[896] = 12'b111111111111;
assign Lowerletter[897] = 12'b111111111111;
assign Lowerletter[898] = 12'b111111111111;
assign Lowerletter[899] = 12'b111111111111;
assign Lowerletter[900] = 12'b111111111111;
assign Lowerletter[901] = 12'b111111111111;
assign Lowerletter[902] = 12'b111111111111;
assign Lowerletter[903] = 12'b111111111111;
assign Lowerletter[904] = 12'b111111111111;
assign Lowerletter[905] = 12'b111111111111;
assign Lowerletter[906] = 12'b111111111111;
assign Lowerletter[907] = 12'b111111111111;
assign Lowerletter[908] = 12'b111111111111;
assign Lowerletter[909] = 12'b111111111111;
assign Lowerletter[910] = 12'b111111111111;
assign Lowerletter[911] = 12'b111111111111;
assign Lowerletter[912] = 12'b111111111111;
assign Lowerletter[913] = 12'b111111111111;
assign Lowerletter[914] = 12'b111111111111;
assign Lowerletter[915] = 12'b000000000000;
assign Lowerletter[916] = 12'b000000000000;
assign Lowerletter[917] = 12'b111111111111;
assign Lowerletter[918] = 12'b111111111111;
assign Lowerletter[919] = 12'b111111111111;
assign Lowerletter[920] = 12'b111111111111;
assign Lowerletter[921] = 12'b111111111111;
assign Lowerletter[922] = 12'b000000000000;
assign Lowerletter[923] = 12'b111111111111;
assign Lowerletter[924] = 12'b111111111111;
assign Lowerletter[925] = 12'b000000000000;
assign Lowerletter[926] = 12'b111111111111;
assign Lowerletter[927] = 12'b111111111111;
assign Lowerletter[928] = 12'b111111111111;
assign Lowerletter[929] = 12'b111111111111;
assign Lowerletter[930] = 12'b000000000000;
assign Lowerletter[931] = 12'b111111111111;
assign Lowerletter[932] = 12'b111111111111;
assign Lowerletter[933] = 12'b000000000000;
assign Lowerletter[934] = 12'b111111111111;
assign Lowerletter[935] = 12'b111111111111;
assign Lowerletter[936] = 12'b111111111111;
assign Lowerletter[937] = 12'b111111111111;
assign Lowerletter[938] = 12'b000000000000;
assign Lowerletter[939] = 12'b111111111111;
assign Lowerletter[940] = 12'b111111111111;
assign Lowerletter[941] = 12'b000000000000;
assign Lowerletter[942] = 12'b111111111111;
assign Lowerletter[943] = 12'b111111111111;
assign Lowerletter[944] = 12'b111111111111;
assign Lowerletter[945] = 12'b111111111111;
assign Lowerletter[946] = 12'b111111111111;
assign Lowerletter[947] = 12'b000000000000;
assign Lowerletter[948] = 12'b000000000000;
assign Lowerletter[949] = 12'b111111111111;
assign Lowerletter[950] = 12'b111111111111;
assign Lowerletter[951] = 12'b111111111111;
assign Lowerletter[952] = 12'b111111111111;
assign Lowerletter[953] = 12'b111111111111;
assign Lowerletter[954] = 12'b111111111111;
assign Lowerletter[955] = 12'b111111111111;
assign Lowerletter[956] = 12'b111111111111;
assign Lowerletter[957] = 12'b111111111111;
assign Lowerletter[958] = 12'b111111111111;
assign Lowerletter[959] = 12'b111111111111;
assign Lowerletter[960] = 12'b111111111111;
assign Lowerletter[961] = 12'b111111111111;
assign Lowerletter[962] = 12'b111111111111;
assign Lowerletter[963] = 12'b111111111111;
assign Lowerletter[964] = 12'b111111111111;
assign Lowerletter[965] = 12'b111111111111;
assign Lowerletter[966] = 12'b111111111111;
assign Lowerletter[967] = 12'b111111111111;
assign Lowerletter[968] = 12'b111111111111;
assign Lowerletter[969] = 12'b111111111111;
assign Lowerletter[970] = 12'b111111111111;
assign Lowerletter[971] = 12'b111111111111;
assign Lowerletter[972] = 12'b111111111111;
assign Lowerletter[973] = 12'b111111111111;
assign Lowerletter[974] = 12'b111111111111;
assign Lowerletter[975] = 12'b111111111111;
assign Lowerletter[976] = 12'b111111111111;
assign Lowerletter[977] = 12'b111111111111;
assign Lowerletter[978] = 12'b000000000000;
assign Lowerletter[979] = 12'b111111111111;
assign Lowerletter[980] = 12'b000000000000;
assign Lowerletter[981] = 12'b111111111111;
assign Lowerletter[982] = 12'b111111111111;
assign Lowerletter[983] = 12'b111111111111;
assign Lowerletter[984] = 12'b111111111111;
assign Lowerletter[985] = 12'b111111111111;
assign Lowerletter[986] = 12'b000000000000;
assign Lowerletter[987] = 12'b000000000000;
assign Lowerletter[988] = 12'b111111111111;
assign Lowerletter[989] = 12'b000000000000;
assign Lowerletter[990] = 12'b111111111111;
assign Lowerletter[991] = 12'b111111111111;
assign Lowerletter[992] = 12'b111111111111;
assign Lowerletter[993] = 12'b111111111111;
assign Lowerletter[994] = 12'b000000000000;
assign Lowerletter[995] = 12'b111111111111;
assign Lowerletter[996] = 12'b111111111111;
assign Lowerletter[997] = 12'b000000000000;
assign Lowerletter[998] = 12'b111111111111;
assign Lowerletter[999] = 12'b111111111111;
assign Lowerletter[1000] = 12'b111111111111;
assign Lowerletter[1001] = 12'b111111111111;
assign Lowerletter[1002] = 12'b000000000000;
assign Lowerletter[1003] = 12'b000000000000;
assign Lowerletter[1004] = 12'b000000000000;
assign Lowerletter[1005] = 12'b111111111111;
assign Lowerletter[1006] = 12'b111111111111;
assign Lowerletter[1007] = 12'b111111111111;
assign Lowerletter[1008] = 12'b111111111111;
assign Lowerletter[1009] = 12'b111111111111;
assign Lowerletter[1010] = 12'b000000000000;
assign Lowerletter[1011] = 12'b111111111111;
assign Lowerletter[1012] = 12'b111111111111;
assign Lowerletter[1013] = 12'b111111111111;
assign Lowerletter[1014] = 12'b111111111111;
assign Lowerletter[1015] = 12'b111111111111;
assign Lowerletter[1016] = 12'b111111111111;
assign Lowerletter[1017] = 12'b111111111111;
assign Lowerletter[1018] = 12'b000000000000;
assign Lowerletter[1019] = 12'b111111111111;
assign Lowerletter[1020] = 12'b111111111111;
assign Lowerletter[1021] = 12'b111111111111;
assign Lowerletter[1022] = 12'b111111111111;
assign Lowerletter[1023] = 12'b111111111111;
assign Lowerletter[1024] = 12'b111111111111;
assign Lowerletter[1025] = 12'b111111111111;
assign Lowerletter[1026] = 12'b111111111111;
assign Lowerletter[1027] = 12'b111111111111;
assign Lowerletter[1028] = 12'b111111111111;
assign Lowerletter[1029] = 12'b111111111111;
assign Lowerletter[1030] = 12'b111111111111;
assign Lowerletter[1031] = 12'b111111111111;
assign Lowerletter[1032] = 12'b111111111111;
assign Lowerletter[1033] = 12'b111111111111;
assign Lowerletter[1034] = 12'b111111111111;
assign Lowerletter[1035] = 12'b111111111111;
assign Lowerletter[1036] = 12'b111111111111;
assign Lowerletter[1037] = 12'b111111111111;
assign Lowerletter[1038] = 12'b111111111111;
assign Lowerletter[1039] = 12'b111111111111;
assign Lowerletter[1040] = 12'b111111111111;
assign Lowerletter[1041] = 12'b111111111111;
assign Lowerletter[1042] = 12'b111111111111;
assign Lowerletter[1043] = 12'b000000000000;
assign Lowerletter[1044] = 12'b111111111111;
assign Lowerletter[1045] = 12'b000000000000;
assign Lowerletter[1046] = 12'b111111111111;
assign Lowerletter[1047] = 12'b111111111111;
assign Lowerletter[1048] = 12'b111111111111;
assign Lowerletter[1049] = 12'b111111111111;
assign Lowerletter[1050] = 12'b000000000000;
assign Lowerletter[1051] = 12'b111111111111;
assign Lowerletter[1052] = 12'b000000000000;
assign Lowerletter[1053] = 12'b000000000000;
assign Lowerletter[1054] = 12'b111111111111;
assign Lowerletter[1055] = 12'b111111111111;
assign Lowerletter[1056] = 12'b111111111111;
assign Lowerletter[1057] = 12'b111111111111;
assign Lowerletter[1058] = 12'b000000000000;
assign Lowerletter[1059] = 12'b111111111111;
assign Lowerletter[1060] = 12'b111111111111;
assign Lowerletter[1061] = 12'b000000000000;
assign Lowerletter[1062] = 12'b111111111111;
assign Lowerletter[1063] = 12'b111111111111;
assign Lowerletter[1064] = 12'b111111111111;
assign Lowerletter[1065] = 12'b111111111111;
assign Lowerletter[1066] = 12'b111111111111;
assign Lowerletter[1067] = 12'b000000000000;
assign Lowerletter[1068] = 12'b000000000000;
assign Lowerletter[1069] = 12'b000000000000;
assign Lowerletter[1070] = 12'b111111111111;
assign Lowerletter[1071] = 12'b111111111111;
assign Lowerletter[1072] = 12'b111111111111;
assign Lowerletter[1073] = 12'b111111111111;
assign Lowerletter[1074] = 12'b111111111111;
assign Lowerletter[1075] = 12'b111111111111;
assign Lowerletter[1076] = 12'b111111111111;
assign Lowerletter[1077] = 12'b000000000000;
assign Lowerletter[1078] = 12'b111111111111;
assign Lowerletter[1079] = 12'b111111111111;
assign Lowerletter[1080] = 12'b111111111111;
assign Lowerletter[1081] = 12'b111111111111;
assign Lowerletter[1082] = 12'b111111111111;
assign Lowerletter[1083] = 12'b111111111111;
assign Lowerletter[1084] = 12'b111111111111;
assign Lowerletter[1085] = 12'b000000000000;
assign Lowerletter[1086] = 12'b111111111111;
assign Lowerletter[1087] = 12'b111111111111;
assign Lowerletter[1088] = 12'b111111111111;
assign Lowerletter[1089] = 12'b111111111111;
assign Lowerletter[1090] = 12'b111111111111;
assign Lowerletter[1091] = 12'b111111111111;
assign Lowerletter[1092] = 12'b111111111111;
assign Lowerletter[1093] = 12'b111111111111;
assign Lowerletter[1094] = 12'b111111111111;
assign Lowerletter[1095] = 12'b111111111111;
assign Lowerletter[1096] = 12'b111111111111;
assign Lowerletter[1097] = 12'b111111111111;
assign Lowerletter[1098] = 12'b111111111111;
assign Lowerletter[1099] = 12'b111111111111;
assign Lowerletter[1100] = 12'b111111111111;
assign Lowerletter[1101] = 12'b111111111111;
assign Lowerletter[1102] = 12'b111111111111;
assign Lowerletter[1103] = 12'b111111111111;
assign Lowerletter[1104] = 12'b111111111111;
assign Lowerletter[1105] = 12'b111111111111;
assign Lowerletter[1106] = 12'b000000000000;
assign Lowerletter[1107] = 12'b111111111111;
assign Lowerletter[1108] = 12'b000000000000;
assign Lowerletter[1109] = 12'b000000000000;
assign Lowerletter[1110] = 12'b111111111111;
assign Lowerletter[1111] = 12'b111111111111;
assign Lowerletter[1112] = 12'b111111111111;
assign Lowerletter[1113] = 12'b111111111111;
assign Lowerletter[1114] = 12'b000000000000;
assign Lowerletter[1115] = 12'b000000000000;
assign Lowerletter[1116] = 12'b111111111111;
assign Lowerletter[1117] = 12'b111111111111;
assign Lowerletter[1118] = 12'b111111111111;
assign Lowerletter[1119] = 12'b111111111111;
assign Lowerletter[1120] = 12'b111111111111;
assign Lowerletter[1121] = 12'b111111111111;
assign Lowerletter[1122] = 12'b000000000000;
assign Lowerletter[1123] = 12'b111111111111;
assign Lowerletter[1124] = 12'b111111111111;
assign Lowerletter[1125] = 12'b111111111111;
assign Lowerletter[1126] = 12'b111111111111;
assign Lowerletter[1127] = 12'b111111111111;
assign Lowerletter[1128] = 12'b111111111111;
assign Lowerletter[1129] = 12'b111111111111;
assign Lowerletter[1130] = 12'b000000000000;
assign Lowerletter[1131] = 12'b111111111111;
assign Lowerletter[1132] = 12'b111111111111;
assign Lowerletter[1133] = 12'b111111111111;
assign Lowerletter[1134] = 12'b111111111111;
assign Lowerletter[1135] = 12'b111111111111;
assign Lowerletter[1136] = 12'b111111111111;
assign Lowerletter[1137] = 12'b111111111111;
assign Lowerletter[1138] = 12'b000000000000;
assign Lowerletter[1139] = 12'b111111111111;
assign Lowerletter[1140] = 12'b111111111111;
assign Lowerletter[1141] = 12'b111111111111;
assign Lowerletter[1142] = 12'b111111111111;
assign Lowerletter[1143] = 12'b111111111111;
assign Lowerletter[1144] = 12'b111111111111;
assign Lowerletter[1145] = 12'b111111111111;
assign Lowerletter[1146] = 12'b111111111111;
assign Lowerletter[1147] = 12'b111111111111;
assign Lowerletter[1148] = 12'b111111111111;
assign Lowerletter[1149] = 12'b111111111111;
assign Lowerletter[1150] = 12'b111111111111;
assign Lowerletter[1151] = 12'b111111111111;
assign Lowerletter[1152] = 12'b111111111111;
assign Lowerletter[1153] = 12'b111111111111;
assign Lowerletter[1154] = 12'b111111111111;
assign Lowerletter[1155] = 12'b111111111111;
assign Lowerletter[1156] = 12'b111111111111;
assign Lowerletter[1157] = 12'b111111111111;
assign Lowerletter[1158] = 12'b111111111111;
assign Lowerletter[1159] = 12'b111111111111;
assign Lowerletter[1160] = 12'b111111111111;
assign Lowerletter[1161] = 12'b111111111111;
assign Lowerletter[1162] = 12'b111111111111;
assign Lowerletter[1163] = 12'b111111111111;
assign Lowerletter[1164] = 12'b111111111111;
assign Lowerletter[1165] = 12'b111111111111;
assign Lowerletter[1166] = 12'b111111111111;
assign Lowerletter[1167] = 12'b111111111111;
assign Lowerletter[1168] = 12'b111111111111;
assign Lowerletter[1169] = 12'b111111111111;
assign Lowerletter[1170] = 12'b111111111111;
assign Lowerletter[1171] = 12'b000000000000;
assign Lowerletter[1172] = 12'b000000000000;
assign Lowerletter[1173] = 12'b000000000000;
assign Lowerletter[1174] = 12'b111111111111;
assign Lowerletter[1175] = 12'b111111111111;
assign Lowerletter[1176] = 12'b111111111111;
assign Lowerletter[1177] = 12'b111111111111;
assign Lowerletter[1178] = 12'b000000000000;
assign Lowerletter[1179] = 12'b111111111111;
assign Lowerletter[1180] = 12'b111111111111;
assign Lowerletter[1181] = 12'b111111111111;
assign Lowerletter[1182] = 12'b111111111111;
assign Lowerletter[1183] = 12'b111111111111;
assign Lowerletter[1184] = 12'b111111111111;
assign Lowerletter[1185] = 12'b111111111111;
assign Lowerletter[1186] = 12'b111111111111;
assign Lowerletter[1187] = 12'b000000000000;
assign Lowerletter[1188] = 12'b000000000000;
assign Lowerletter[1189] = 12'b111111111111;
assign Lowerletter[1190] = 12'b111111111111;
assign Lowerletter[1191] = 12'b111111111111;
assign Lowerletter[1192] = 12'b111111111111;
assign Lowerletter[1193] = 12'b111111111111;
assign Lowerletter[1194] = 12'b111111111111;
assign Lowerletter[1195] = 12'b111111111111;
assign Lowerletter[1196] = 12'b111111111111;
assign Lowerletter[1197] = 12'b000000000000;
assign Lowerletter[1198] = 12'b111111111111;
assign Lowerletter[1199] = 12'b111111111111;
assign Lowerletter[1200] = 12'b111111111111;
assign Lowerletter[1201] = 12'b111111111111;
assign Lowerletter[1202] = 12'b000000000000;
assign Lowerletter[1203] = 12'b000000000000;
assign Lowerletter[1204] = 12'b000000000000;
assign Lowerletter[1205] = 12'b111111111111;
assign Lowerletter[1206] = 12'b111111111111;
assign Lowerletter[1207] = 12'b111111111111;
assign Lowerletter[1208] = 12'b111111111111;
assign Lowerletter[1209] = 12'b111111111111;
assign Lowerletter[1210] = 12'b111111111111;
assign Lowerletter[1211] = 12'b111111111111;
assign Lowerletter[1212] = 12'b111111111111;
assign Lowerletter[1213] = 12'b111111111111;
assign Lowerletter[1214] = 12'b111111111111;
assign Lowerletter[1215] = 12'b111111111111;
assign Lowerletter[1216] = 12'b111111111111;
assign Lowerletter[1217] = 12'b111111111111;
assign Lowerletter[1218] = 12'b111111111111;
assign Lowerletter[1219] = 12'b111111111111;
assign Lowerletter[1220] = 12'b111111111111;
assign Lowerletter[1221] = 12'b111111111111;
assign Lowerletter[1222] = 12'b111111111111;
assign Lowerletter[1223] = 12'b111111111111;
assign Lowerletter[1224] = 12'b111111111111;
assign Lowerletter[1225] = 12'b111111111111;
assign Lowerletter[1226] = 12'b111111111111;
assign Lowerletter[1227] = 12'b000000000000;
assign Lowerletter[1228] = 12'b111111111111;
assign Lowerletter[1229] = 12'b111111111111;
assign Lowerletter[1230] = 12'b111111111111;
assign Lowerletter[1231] = 12'b111111111111;
assign Lowerletter[1232] = 12'b111111111111;
assign Lowerletter[1233] = 12'b111111111111;
assign Lowerletter[1234] = 12'b000000000000;
assign Lowerletter[1235] = 12'b000000000000;
assign Lowerletter[1236] = 12'b000000000000;
assign Lowerletter[1237] = 12'b111111111111;
assign Lowerletter[1238] = 12'b111111111111;
assign Lowerletter[1239] = 12'b111111111111;
assign Lowerletter[1240] = 12'b111111111111;
assign Lowerletter[1241] = 12'b111111111111;
assign Lowerletter[1242] = 12'b111111111111;
assign Lowerletter[1243] = 12'b000000000000;
assign Lowerletter[1244] = 12'b111111111111;
assign Lowerletter[1245] = 12'b111111111111;
assign Lowerletter[1246] = 12'b111111111111;
assign Lowerletter[1247] = 12'b111111111111;
assign Lowerletter[1248] = 12'b111111111111;
assign Lowerletter[1249] = 12'b111111111111;
assign Lowerletter[1250] = 12'b111111111111;
assign Lowerletter[1251] = 12'b000000000000;
assign Lowerletter[1252] = 12'b111111111111;
assign Lowerletter[1253] = 12'b111111111111;
assign Lowerletter[1254] = 12'b111111111111;
assign Lowerletter[1255] = 12'b111111111111;
assign Lowerletter[1256] = 12'b111111111111;
assign Lowerletter[1257] = 12'b111111111111;
assign Lowerletter[1258] = 12'b111111111111;
assign Lowerletter[1259] = 12'b000000000000;
assign Lowerletter[1260] = 12'b111111111111;
assign Lowerletter[1261] = 12'b111111111111;
assign Lowerletter[1262] = 12'b111111111111;
assign Lowerletter[1263] = 12'b111111111111;
assign Lowerletter[1264] = 12'b111111111111;
assign Lowerletter[1265] = 12'b111111111111;
assign Lowerletter[1266] = 12'b111111111111;
assign Lowerletter[1267] = 12'b111111111111;
assign Lowerletter[1268] = 12'b000000000000;
assign Lowerletter[1269] = 12'b111111111111;
assign Lowerletter[1270] = 12'b111111111111;
assign Lowerletter[1271] = 12'b111111111111;
assign Lowerletter[1272] = 12'b111111111111;
assign Lowerletter[1273] = 12'b111111111111;
assign Lowerletter[1274] = 12'b111111111111;
assign Lowerletter[1275] = 12'b111111111111;
assign Lowerletter[1276] = 12'b111111111111;
assign Lowerletter[1277] = 12'b111111111111;
assign Lowerletter[1278] = 12'b111111111111;
assign Lowerletter[1279] = 12'b111111111111;
assign Lowerletter[1280] = 12'b111111111111;
assign Lowerletter[1281] = 12'b111111111111;
assign Lowerletter[1282] = 12'b111111111111;
assign Lowerletter[1283] = 12'b111111111111;
assign Lowerletter[1284] = 12'b111111111111;
assign Lowerletter[1285] = 12'b111111111111;
assign Lowerletter[1286] = 12'b111111111111;
assign Lowerletter[1287] = 12'b111111111111;
assign Lowerletter[1288] = 12'b111111111111;
assign Lowerletter[1289] = 12'b111111111111;
assign Lowerletter[1290] = 12'b111111111111;
assign Lowerletter[1291] = 12'b111111111111;
assign Lowerletter[1292] = 12'b111111111111;
assign Lowerletter[1293] = 12'b111111111111;
assign Lowerletter[1294] = 12'b111111111111;
assign Lowerletter[1295] = 12'b111111111111;
assign Lowerletter[1296] = 12'b111111111111;
assign Lowerletter[1297] = 12'b111111111111;
assign Lowerletter[1298] = 12'b000000000000;
assign Lowerletter[1299] = 12'b111111111111;
assign Lowerletter[1300] = 12'b111111111111;
assign Lowerletter[1301] = 12'b000000000000;
assign Lowerletter[1302] = 12'b111111111111;
assign Lowerletter[1303] = 12'b111111111111;
assign Lowerletter[1304] = 12'b111111111111;
assign Lowerletter[1305] = 12'b111111111111;
assign Lowerletter[1306] = 12'b000000000000;
assign Lowerletter[1307] = 12'b111111111111;
assign Lowerletter[1308] = 12'b111111111111;
assign Lowerletter[1309] = 12'b000000000000;
assign Lowerletter[1310] = 12'b111111111111;
assign Lowerletter[1311] = 12'b111111111111;
assign Lowerletter[1312] = 12'b111111111111;
assign Lowerletter[1313] = 12'b111111111111;
assign Lowerletter[1314] = 12'b000000000000;
assign Lowerletter[1315] = 12'b111111111111;
assign Lowerletter[1316] = 12'b111111111111;
assign Lowerletter[1317] = 12'b000000000000;
assign Lowerletter[1318] = 12'b111111111111;
assign Lowerletter[1319] = 12'b111111111111;
assign Lowerletter[1320] = 12'b111111111111;
assign Lowerletter[1321] = 12'b111111111111;
assign Lowerletter[1322] = 12'b000000000000;
assign Lowerletter[1323] = 12'b111111111111;
assign Lowerletter[1324] = 12'b111111111111;
assign Lowerletter[1325] = 12'b000000000000;
assign Lowerletter[1326] = 12'b111111111111;
assign Lowerletter[1327] = 12'b111111111111;
assign Lowerletter[1328] = 12'b111111111111;
assign Lowerletter[1329] = 12'b111111111111;
assign Lowerletter[1330] = 12'b111111111111;
assign Lowerletter[1331] = 12'b000000000000;
assign Lowerletter[1332] = 12'b000000000000;
assign Lowerletter[1333] = 12'b111111111111;
assign Lowerletter[1334] = 12'b111111111111;
assign Lowerletter[1335] = 12'b111111111111;
assign Lowerletter[1336] = 12'b111111111111;
assign Lowerletter[1337] = 12'b111111111111;
assign Lowerletter[1338] = 12'b111111111111;
assign Lowerletter[1339] = 12'b111111111111;
assign Lowerletter[1340] = 12'b111111111111;
assign Lowerletter[1341] = 12'b111111111111;
assign Lowerletter[1342] = 12'b111111111111;
assign Lowerletter[1343] = 12'b111111111111;
assign Lowerletter[1344] = 12'b111111111111;
assign Lowerletter[1345] = 12'b111111111111;
assign Lowerletter[1346] = 12'b111111111111;
assign Lowerletter[1347] = 12'b111111111111;
assign Lowerletter[1348] = 12'b111111111111;
assign Lowerletter[1349] = 12'b111111111111;
assign Lowerletter[1350] = 12'b111111111111;
assign Lowerletter[1351] = 12'b111111111111;
assign Lowerletter[1352] = 12'b111111111111;
assign Lowerletter[1353] = 12'b111111111111;
assign Lowerletter[1354] = 12'b111111111111;
assign Lowerletter[1355] = 12'b111111111111;
assign Lowerletter[1356] = 12'b111111111111;
assign Lowerletter[1357] = 12'b111111111111;
assign Lowerletter[1358] = 12'b111111111111;
assign Lowerletter[1359] = 12'b111111111111;
assign Lowerletter[1360] = 12'b111111111111;
assign Lowerletter[1361] = 12'b000000000000;
assign Lowerletter[1362] = 12'b111111111111;
assign Lowerletter[1363] = 12'b111111111111;
assign Lowerletter[1364] = 12'b111111111111;
assign Lowerletter[1365] = 12'b000000000000;
assign Lowerletter[1366] = 12'b111111111111;
assign Lowerletter[1367] = 12'b111111111111;
assign Lowerletter[1368] = 12'b111111111111;
assign Lowerletter[1369] = 12'b000000000000;
assign Lowerletter[1370] = 12'b111111111111;
assign Lowerletter[1371] = 12'b111111111111;
assign Lowerletter[1372] = 12'b111111111111;
assign Lowerletter[1373] = 12'b000000000000;
assign Lowerletter[1374] = 12'b111111111111;
assign Lowerletter[1375] = 12'b111111111111;
assign Lowerletter[1376] = 12'b111111111111;
assign Lowerletter[1377] = 12'b000000000000;
assign Lowerletter[1378] = 12'b111111111111;
assign Lowerletter[1379] = 12'b111111111111;
assign Lowerletter[1380] = 12'b111111111111;
assign Lowerletter[1381] = 12'b000000000000;
assign Lowerletter[1382] = 12'b111111111111;
assign Lowerletter[1383] = 12'b111111111111;
assign Lowerletter[1384] = 12'b111111111111;
assign Lowerletter[1385] = 12'b111111111111;
assign Lowerletter[1386] = 12'b000000000000;
assign Lowerletter[1387] = 12'b111111111111;
assign Lowerletter[1388] = 12'b000000000000;
assign Lowerletter[1389] = 12'b111111111111;
assign Lowerletter[1390] = 12'b111111111111;
assign Lowerletter[1391] = 12'b111111111111;
assign Lowerletter[1392] = 12'b111111111111;
assign Lowerletter[1393] = 12'b111111111111;
assign Lowerletter[1394] = 12'b111111111111;
assign Lowerletter[1395] = 12'b000000000000;
assign Lowerletter[1396] = 12'b111111111111;
assign Lowerletter[1397] = 12'b111111111111;
assign Lowerletter[1398] = 12'b111111111111;
assign Lowerletter[1399] = 12'b111111111111;
assign Lowerletter[1400] = 12'b111111111111;
assign Lowerletter[1401] = 12'b111111111111;
assign Lowerletter[1402] = 12'b111111111111;
assign Lowerletter[1403] = 12'b111111111111;
assign Lowerletter[1404] = 12'b111111111111;
assign Lowerletter[1405] = 12'b111111111111;
assign Lowerletter[1406] = 12'b111111111111;
assign Lowerletter[1407] = 12'b111111111111;
assign Lowerletter[1408] = 12'b111111111111;
assign Lowerletter[1409] = 12'b111111111111;
assign Lowerletter[1410] = 12'b111111111111;
assign Lowerletter[1411] = 12'b111111111111;
assign Lowerletter[1412] = 12'b111111111111;
assign Lowerletter[1413] = 12'b111111111111;
assign Lowerletter[1414] = 12'b111111111111;
assign Lowerletter[1415] = 12'b111111111111;
assign Lowerletter[1416] = 12'b111111111111;
assign Lowerletter[1417] = 12'b111111111111;
assign Lowerletter[1418] = 12'b111111111111;
assign Lowerletter[1419] = 12'b111111111111;
assign Lowerletter[1420] = 12'b111111111111;
assign Lowerletter[1421] = 12'b111111111111;
assign Lowerletter[1422] = 12'b111111111111;
assign Lowerletter[1423] = 12'b111111111111;
assign Lowerletter[1424] = 12'b111111111111;
assign Lowerletter[1425] = 12'b111111111111;
assign Lowerletter[1426] = 12'b111111111111;
assign Lowerletter[1427] = 12'b111111111111;
assign Lowerletter[1428] = 12'b111111111111;
assign Lowerletter[1429] = 12'b111111111111;
assign Lowerletter[1430] = 12'b111111111111;
assign Lowerletter[1431] = 12'b111111111111;
assign Lowerletter[1432] = 12'b111111111111;
assign Lowerletter[1433] = 12'b000000000000;
assign Lowerletter[1434] = 12'b111111111111;
assign Lowerletter[1435] = 12'b111111111111;
assign Lowerletter[1436] = 12'b111111111111;
assign Lowerletter[1437] = 12'b000000000000;
assign Lowerletter[1438] = 12'b111111111111;
assign Lowerletter[1439] = 12'b111111111111;
assign Lowerletter[1440] = 12'b111111111111;
assign Lowerletter[1441] = 12'b000000000000;
assign Lowerletter[1442] = 12'b111111111111;
assign Lowerletter[1443] = 12'b111111111111;
assign Lowerletter[1444] = 12'b111111111111;
assign Lowerletter[1445] = 12'b000000000000;
assign Lowerletter[1446] = 12'b111111111111;
assign Lowerletter[1447] = 12'b111111111111;
assign Lowerletter[1448] = 12'b111111111111;
assign Lowerletter[1449] = 12'b000000000000;
assign Lowerletter[1450] = 12'b111111111111;
assign Lowerletter[1451] = 12'b000000000000;
assign Lowerletter[1452] = 12'b111111111111;
assign Lowerletter[1453] = 12'b000000000000;
assign Lowerletter[1454] = 12'b111111111111;
assign Lowerletter[1455] = 12'b111111111111;
assign Lowerletter[1456] = 12'b111111111111;
assign Lowerletter[1457] = 12'b111111111111;
assign Lowerletter[1458] = 12'b000000000000;
assign Lowerletter[1459] = 12'b000000000000;
assign Lowerletter[1460] = 12'b000000000000;
assign Lowerletter[1461] = 12'b000000000000;
assign Lowerletter[1462] = 12'b111111111111;
assign Lowerletter[1463] = 12'b111111111111;
assign Lowerletter[1464] = 12'b111111111111;
assign Lowerletter[1465] = 12'b111111111111;
assign Lowerletter[1466] = 12'b111111111111;
assign Lowerletter[1467] = 12'b111111111111;
assign Lowerletter[1468] = 12'b111111111111;
assign Lowerletter[1469] = 12'b111111111111;
assign Lowerletter[1470] = 12'b111111111111;
assign Lowerletter[1471] = 12'b111111111111;
assign Lowerletter[1472] = 12'b111111111111;
assign Lowerletter[1473] = 12'b111111111111;
assign Lowerletter[1474] = 12'b111111111111;
assign Lowerletter[1475] = 12'b111111111111;
assign Lowerletter[1476] = 12'b111111111111;
assign Lowerletter[1477] = 12'b111111111111;
assign Lowerletter[1478] = 12'b111111111111;
assign Lowerletter[1479] = 12'b111111111111;
assign Lowerletter[1480] = 12'b111111111111;
assign Lowerletter[1481] = 12'b111111111111;
assign Lowerletter[1482] = 12'b111111111111;
assign Lowerletter[1483] = 12'b111111111111;
assign Lowerletter[1484] = 12'b111111111111;
assign Lowerletter[1485] = 12'b111111111111;
assign Lowerletter[1486] = 12'b111111111111;
assign Lowerletter[1487] = 12'b111111111111;
assign Lowerletter[1488] = 12'b111111111111;
assign Lowerletter[1489] = 12'b000000000000;
assign Lowerletter[1490] = 12'b111111111111;
assign Lowerletter[1491] = 12'b111111111111;
assign Lowerletter[1492] = 12'b111111111111;
assign Lowerletter[1493] = 12'b000000000000;
assign Lowerletter[1494] = 12'b111111111111;
assign Lowerletter[1495] = 12'b111111111111;
assign Lowerletter[1496] = 12'b111111111111;
assign Lowerletter[1497] = 12'b111111111111;
assign Lowerletter[1498] = 12'b000000000000;
assign Lowerletter[1499] = 12'b111111111111;
assign Lowerletter[1500] = 12'b000000000000;
assign Lowerletter[1501] = 12'b111111111111;
assign Lowerletter[1502] = 12'b111111111111;
assign Lowerletter[1503] = 12'b111111111111;
assign Lowerletter[1504] = 12'b111111111111;
assign Lowerletter[1505] = 12'b111111111111;
assign Lowerletter[1506] = 12'b111111111111;
assign Lowerletter[1507] = 12'b000000000000;
assign Lowerletter[1508] = 12'b111111111111;
assign Lowerletter[1509] = 12'b111111111111;
assign Lowerletter[1510] = 12'b111111111111;
assign Lowerletter[1511] = 12'b111111111111;
assign Lowerletter[1512] = 12'b111111111111;
assign Lowerletter[1513] = 12'b111111111111;
assign Lowerletter[1514] = 12'b000000000000;
assign Lowerletter[1515] = 12'b111111111111;
assign Lowerletter[1516] = 12'b000000000000;
assign Lowerletter[1517] = 12'b111111111111;
assign Lowerletter[1518] = 12'b111111111111;
assign Lowerletter[1519] = 12'b111111111111;
assign Lowerletter[1520] = 12'b111111111111;
assign Lowerletter[1521] = 12'b000000000000;
assign Lowerletter[1522] = 12'b111111111111;
assign Lowerletter[1523] = 12'b111111111111;
assign Lowerletter[1524] = 12'b111111111111;
assign Lowerletter[1525] = 12'b000000000000;
assign Lowerletter[1526] = 12'b111111111111;
assign Lowerletter[1527] = 12'b111111111111;
assign Lowerletter[1528] = 12'b111111111111;
assign Lowerletter[1529] = 12'b111111111111;
assign Lowerletter[1530] = 12'b111111111111;
assign Lowerletter[1531] = 12'b111111111111;
assign Lowerletter[1532] = 12'b111111111111;
assign Lowerletter[1533] = 12'b111111111111;
assign Lowerletter[1534] = 12'b111111111111;
assign Lowerletter[1535] = 12'b111111111111;
assign Lowerletter[1536] = 12'b111111111111;
assign Lowerletter[1537] = 12'b111111111111;
assign Lowerletter[1538] = 12'b111111111111;
assign Lowerletter[1539] = 12'b111111111111;
assign Lowerletter[1540] = 12'b111111111111;
assign Lowerletter[1541] = 12'b111111111111;
assign Lowerletter[1542] = 12'b111111111111;
assign Lowerletter[1543] = 12'b111111111111;
assign Lowerletter[1544] = 12'b111111111111;
assign Lowerletter[1545] = 12'b111111111111;
assign Lowerletter[1546] = 12'b111111111111;
assign Lowerletter[1547] = 12'b111111111111;
assign Lowerletter[1548] = 12'b111111111111;
assign Lowerletter[1549] = 12'b111111111111;
assign Lowerletter[1550] = 12'b111111111111;
assign Lowerletter[1551] = 12'b111111111111;
assign Lowerletter[1552] = 12'b111111111111;
assign Lowerletter[1553] = 12'b111111111111;
assign Lowerletter[1554] = 12'b000000000000;
assign Lowerletter[1555] = 12'b111111111111;
assign Lowerletter[1556] = 12'b111111111111;
assign Lowerletter[1557] = 12'b000000000000;
assign Lowerletter[1558] = 12'b111111111111;
assign Lowerletter[1559] = 12'b111111111111;
assign Lowerletter[1560] = 12'b111111111111;
assign Lowerletter[1561] = 12'b111111111111;
assign Lowerletter[1562] = 12'b000000000000;
assign Lowerletter[1563] = 12'b111111111111;
assign Lowerletter[1564] = 12'b111111111111;
assign Lowerletter[1565] = 12'b000000000000;
assign Lowerletter[1566] = 12'b111111111111;
assign Lowerletter[1567] = 12'b111111111111;
assign Lowerletter[1568] = 12'b111111111111;
assign Lowerletter[1569] = 12'b111111111111;
assign Lowerletter[1570] = 12'b000000000000;
assign Lowerletter[1571] = 12'b111111111111;
assign Lowerletter[1572] = 12'b111111111111;
assign Lowerletter[1573] = 12'b000000000000;
assign Lowerletter[1574] = 12'b111111111111;
assign Lowerletter[1575] = 12'b111111111111;
assign Lowerletter[1576] = 12'b111111111111;
assign Lowerletter[1577] = 12'b111111111111;
assign Lowerletter[1578] = 12'b111111111111;
assign Lowerletter[1579] = 12'b000000000000;
assign Lowerletter[1580] = 12'b000000000000;
assign Lowerletter[1581] = 12'b000000000000;
assign Lowerletter[1582] = 12'b111111111111;
assign Lowerletter[1583] = 12'b111111111111;
assign Lowerletter[1584] = 12'b111111111111;
assign Lowerletter[1585] = 12'b111111111111;
assign Lowerletter[1586] = 12'b111111111111;
assign Lowerletter[1587] = 12'b111111111111;
assign Lowerletter[1588] = 12'b111111111111;
assign Lowerletter[1589] = 12'b000000000000;
assign Lowerletter[1590] = 12'b111111111111;
assign Lowerletter[1591] = 12'b111111111111;
assign Lowerletter[1592] = 12'b111111111111;
assign Lowerletter[1593] = 12'b111111111111;
assign Lowerletter[1594] = 12'b000000000000;
assign Lowerletter[1595] = 12'b000000000000;
assign Lowerletter[1596] = 12'b000000000000;
assign Lowerletter[1597] = 12'b111111111111;
assign Lowerletter[1598] = 12'b111111111111;
assign Lowerletter[1599] = 12'b111111111111;
assign Lowerletter[1600] = 12'b111111111111;
assign Lowerletter[1601] = 12'b111111111111;
assign Lowerletter[1602] = 12'b111111111111;
assign Lowerletter[1603] = 12'b111111111111;
assign Lowerletter[1604] = 12'b111111111111;
assign Lowerletter[1605] = 12'b111111111111;
assign Lowerletter[1606] = 12'b111111111111;
assign Lowerletter[1607] = 12'b111111111111;
assign Lowerletter[1608] = 12'b111111111111;
assign Lowerletter[1609] = 12'b111111111111;
assign Lowerletter[1610] = 12'b111111111111;
assign Lowerletter[1611] = 12'b111111111111;
assign Lowerletter[1612] = 12'b111111111111;
assign Lowerletter[1613] = 12'b111111111111;
assign Lowerletter[1614] = 12'b111111111111;
assign Lowerletter[1615] = 12'b111111111111;
assign Lowerletter[1616] = 12'b111111111111;
assign Lowerletter[1617] = 12'b000000000000;
assign Lowerletter[1618] = 12'b000000000000;
assign Lowerletter[1619] = 12'b000000000000;
assign Lowerletter[1620] = 12'b000000000000;
assign Lowerletter[1621] = 12'b000000000000;
assign Lowerletter[1622] = 12'b111111111111;
assign Lowerletter[1623] = 12'b111111111111;
assign Lowerletter[1624] = 12'b111111111111;
assign Lowerletter[1625] = 12'b111111111111;
assign Lowerletter[1626] = 12'b111111111111;
assign Lowerletter[1627] = 12'b111111111111;
assign Lowerletter[1628] = 12'b000000000000;
assign Lowerletter[1629] = 12'b111111111111;
assign Lowerletter[1630] = 12'b111111111111;
assign Lowerletter[1631] = 12'b111111111111;
assign Lowerletter[1632] = 12'b111111111111;
assign Lowerletter[1633] = 12'b111111111111;
assign Lowerletter[1634] = 12'b111111111111;
assign Lowerletter[1635] = 12'b000000000000;
assign Lowerletter[1636] = 12'b111111111111;
assign Lowerletter[1637] = 12'b111111111111;
assign Lowerletter[1638] = 12'b111111111111;
assign Lowerletter[1639] = 12'b111111111111;
assign Lowerletter[1640] = 12'b111111111111;
assign Lowerletter[1641] = 12'b111111111111;
assign Lowerletter[1642] = 12'b000000000000;
assign Lowerletter[1643] = 12'b111111111111;
assign Lowerletter[1644] = 12'b111111111111;
assign Lowerletter[1645] = 12'b111111111111;
assign Lowerletter[1646] = 12'b111111111111;
assign Lowerletter[1647] = 12'b111111111111;
assign Lowerletter[1648] = 12'b111111111111;
assign Lowerletter[1649] = 12'b000000000000;
assign Lowerletter[1650] = 12'b000000000000;
assign Lowerletter[1651] = 12'b000000000000;
assign Lowerletter[1652] = 12'b000000000000;
assign Lowerletter[1653] = 12'b000000000000;
assign Lowerletter[1654] = 12'b111111111111;
assign Lowerletter[1655] = 12'b111111111111;
assign Lowerletter[1656] = 12'b111111111111;
assign Lowerletter[1657] = 12'b111111111111;
assign Lowerletter[1658] = 12'b111111111111;
assign Lowerletter[1659] = 12'b111111111111;
assign Lowerletter[1660] = 12'b111111111111;
assign Lowerletter[1661] = 12'b111111111111;
assign Lowerletter[1662] = 12'b111111111111;
assign Lowerletter[1663] = 12'b111111111111;
assign Upperletter[0] = 12'b111111111111;
assign Upperletter[1] = 12'b111111111111;
assign Upperletter[2] = 12'b000000000000;
assign Upperletter[3] = 12'b000000000000;
assign Upperletter[4] = 12'b000000000000;
assign Upperletter[5] = 12'b111111111111;
assign Upperletter[6] = 12'b111111111111;
assign Upperletter[7] = 12'b111111111111;
assign Upperletter[8] = 12'b111111111111;
assign Upperletter[9] = 12'b000000000000;
assign Upperletter[10] = 12'b111111111111;
assign Upperletter[11] = 12'b111111111111;
assign Upperletter[12] = 12'b111111111111;
assign Upperletter[13] = 12'b000000000000;
assign Upperletter[14] = 12'b111111111111;
assign Upperletter[15] = 12'b111111111111;
assign Upperletter[16] = 12'b111111111111;
assign Upperletter[17] = 12'b000000000000;
assign Upperletter[18] = 12'b111111111111;
assign Upperletter[19] = 12'b111111111111;
assign Upperletter[20] = 12'b111111111111;
assign Upperletter[21] = 12'b000000000000;
assign Upperletter[22] = 12'b111111111111;
assign Upperletter[23] = 12'b111111111111;
assign Upperletter[24] = 12'b111111111111;
assign Upperletter[25] = 12'b000000000000;
assign Upperletter[26] = 12'b000000000000;
assign Upperletter[27] = 12'b000000000000;
assign Upperletter[28] = 12'b000000000000;
assign Upperletter[29] = 12'b000000000000;
assign Upperletter[30] = 12'b111111111111;
assign Upperletter[31] = 12'b111111111111;
assign Upperletter[32] = 12'b111111111111;
assign Upperletter[33] = 12'b000000000000;
assign Upperletter[34] = 12'b111111111111;
assign Upperletter[35] = 12'b111111111111;
assign Upperletter[36] = 12'b111111111111;
assign Upperletter[37] = 12'b000000000000;
assign Upperletter[38] = 12'b111111111111;
assign Upperletter[39] = 12'b111111111111;
assign Upperletter[40] = 12'b111111111111;
assign Upperletter[41] = 12'b000000000000;
assign Upperletter[42] = 12'b111111111111;
assign Upperletter[43] = 12'b111111111111;
assign Upperletter[44] = 12'b111111111111;
assign Upperletter[45] = 12'b000000000000;
assign Upperletter[46] = 12'b111111111111;
assign Upperletter[47] = 12'b111111111111;
assign Upperletter[48] = 12'b111111111111;
assign Upperletter[49] = 12'b000000000000;
assign Upperletter[50] = 12'b111111111111;
assign Upperletter[51] = 12'b111111111111;
assign Upperletter[52] = 12'b111111111111;
assign Upperletter[53] = 12'b000000000000;
assign Upperletter[54] = 12'b111111111111;
assign Upperletter[55] = 12'b111111111111;
assign Upperletter[56] = 12'b111111111111;
assign Upperletter[57] = 12'b111111111111;
assign Upperletter[58] = 12'b111111111111;
assign Upperletter[59] = 12'b111111111111;
assign Upperletter[60] = 12'b111111111111;
assign Upperletter[61] = 12'b111111111111;
assign Upperletter[62] = 12'b111111111111;
assign Upperletter[63] = 12'b111111111111;
assign Upperletter[64] = 12'b111111111111;
assign Upperletter[65] = 12'b000000000000;
assign Upperletter[66] = 12'b000000000000;
assign Upperletter[67] = 12'b000000000000;
assign Upperletter[68] = 12'b000000000000;
assign Upperletter[69] = 12'b111111111111;
assign Upperletter[70] = 12'b111111111111;
assign Upperletter[71] = 12'b111111111111;
assign Upperletter[72] = 12'b111111111111;
assign Upperletter[73] = 12'b000000000000;
assign Upperletter[74] = 12'b111111111111;
assign Upperletter[75] = 12'b111111111111;
assign Upperletter[76] = 12'b111111111111;
assign Upperletter[77] = 12'b000000000000;
assign Upperletter[78] = 12'b111111111111;
assign Upperletter[79] = 12'b111111111111;
assign Upperletter[80] = 12'b111111111111;
assign Upperletter[81] = 12'b000000000000;
assign Upperletter[82] = 12'b111111111111;
assign Upperletter[83] = 12'b111111111111;
assign Upperletter[84] = 12'b111111111111;
assign Upperletter[85] = 12'b000000000000;
assign Upperletter[86] = 12'b111111111111;
assign Upperletter[87] = 12'b111111111111;
assign Upperletter[88] = 12'b111111111111;
assign Upperletter[89] = 12'b000000000000;
assign Upperletter[90] = 12'b000000000000;
assign Upperletter[91] = 12'b000000000000;
assign Upperletter[92] = 12'b000000000000;
assign Upperletter[93] = 12'b111111111111;
assign Upperletter[94] = 12'b111111111111;
assign Upperletter[95] = 12'b111111111111;
assign Upperletter[96] = 12'b111111111111;
assign Upperletter[97] = 12'b000000000000;
assign Upperletter[98] = 12'b111111111111;
assign Upperletter[99] = 12'b111111111111;
assign Upperletter[100] = 12'b111111111111;
assign Upperletter[101] = 12'b000000000000;
assign Upperletter[102] = 12'b111111111111;
assign Upperletter[103] = 12'b111111111111;
assign Upperletter[104] = 12'b111111111111;
assign Upperletter[105] = 12'b000000000000;
assign Upperletter[106] = 12'b111111111111;
assign Upperletter[107] = 12'b111111111111;
assign Upperletter[108] = 12'b111111111111;
assign Upperletter[109] = 12'b000000000000;
assign Upperletter[110] = 12'b111111111111;
assign Upperletter[111] = 12'b111111111111;
assign Upperletter[112] = 12'b111111111111;
assign Upperletter[113] = 12'b000000000000;
assign Upperletter[114] = 12'b000000000000;
assign Upperletter[115] = 12'b000000000000;
assign Upperletter[116] = 12'b000000000000;
assign Upperletter[117] = 12'b111111111111;
assign Upperletter[118] = 12'b111111111111;
assign Upperletter[119] = 12'b111111111111;
assign Upperletter[120] = 12'b111111111111;
assign Upperletter[121] = 12'b111111111111;
assign Upperletter[122] = 12'b111111111111;
assign Upperletter[123] = 12'b111111111111;
assign Upperletter[124] = 12'b111111111111;
assign Upperletter[125] = 12'b111111111111;
assign Upperletter[126] = 12'b111111111111;
assign Upperletter[127] = 12'b111111111111;
assign Upperletter[128] = 12'b111111111111;
assign Upperletter[129] = 12'b111111111111;
assign Upperletter[130] = 12'b000000000000;
assign Upperletter[131] = 12'b000000000000;
assign Upperletter[132] = 12'b000000000000;
assign Upperletter[133] = 12'b111111111111;
assign Upperletter[134] = 12'b111111111111;
assign Upperletter[135] = 12'b111111111111;
assign Upperletter[136] = 12'b111111111111;
assign Upperletter[137] = 12'b000000000000;
assign Upperletter[138] = 12'b111111111111;
assign Upperletter[139] = 12'b111111111111;
assign Upperletter[140] = 12'b111111111111;
assign Upperletter[141] = 12'b000000000000;
assign Upperletter[142] = 12'b111111111111;
assign Upperletter[143] = 12'b111111111111;
assign Upperletter[144] = 12'b111111111111;
assign Upperletter[145] = 12'b000000000000;
assign Upperletter[146] = 12'b111111111111;
assign Upperletter[147] = 12'b111111111111;
assign Upperletter[148] = 12'b111111111111;
assign Upperletter[149] = 12'b111111111111;
assign Upperletter[150] = 12'b111111111111;
assign Upperletter[151] = 12'b111111111111;
assign Upperletter[152] = 12'b111111111111;
assign Upperletter[153] = 12'b000000000000;
assign Upperletter[154] = 12'b111111111111;
assign Upperletter[155] = 12'b111111111111;
assign Upperletter[156] = 12'b111111111111;
assign Upperletter[157] = 12'b111111111111;
assign Upperletter[158] = 12'b111111111111;
assign Upperletter[159] = 12'b111111111111;
assign Upperletter[160] = 12'b111111111111;
assign Upperletter[161] = 12'b000000000000;
assign Upperletter[162] = 12'b111111111111;
assign Upperletter[163] = 12'b111111111111;
assign Upperletter[164] = 12'b111111111111;
assign Upperletter[165] = 12'b111111111111;
assign Upperletter[166] = 12'b111111111111;
assign Upperletter[167] = 12'b111111111111;
assign Upperletter[168] = 12'b111111111111;
assign Upperletter[169] = 12'b000000000000;
assign Upperletter[170] = 12'b111111111111;
assign Upperletter[171] = 12'b111111111111;
assign Upperletter[172] = 12'b111111111111;
assign Upperletter[173] = 12'b000000000000;
assign Upperletter[174] = 12'b111111111111;
assign Upperletter[175] = 12'b111111111111;
assign Upperletter[176] = 12'b111111111111;
assign Upperletter[177] = 12'b111111111111;
assign Upperletter[178] = 12'b000000000000;
assign Upperletter[179] = 12'b000000000000;
assign Upperletter[180] = 12'b000000000000;
assign Upperletter[181] = 12'b111111111111;
assign Upperletter[182] = 12'b111111111111;
assign Upperletter[183] = 12'b111111111111;
assign Upperletter[184] = 12'b111111111111;
assign Upperletter[185] = 12'b111111111111;
assign Upperletter[186] = 12'b111111111111;
assign Upperletter[187] = 12'b111111111111;
assign Upperletter[188] = 12'b111111111111;
assign Upperletter[189] = 12'b111111111111;
assign Upperletter[190] = 12'b111111111111;
assign Upperletter[191] = 12'b111111111111;
assign Upperletter[192] = 12'b111111111111;
assign Upperletter[193] = 12'b000000000000;
assign Upperletter[194] = 12'b000000000000;
assign Upperletter[195] = 12'b000000000000;
assign Upperletter[196] = 12'b000000000000;
assign Upperletter[197] = 12'b111111111111;
assign Upperletter[198] = 12'b111111111111;
assign Upperletter[199] = 12'b111111111111;
assign Upperletter[200] = 12'b111111111111;
assign Upperletter[201] = 12'b000000000000;
assign Upperletter[202] = 12'b111111111111;
assign Upperletter[203] = 12'b111111111111;
assign Upperletter[204] = 12'b111111111111;
assign Upperletter[205] = 12'b000000000000;
assign Upperletter[206] = 12'b111111111111;
assign Upperletter[207] = 12'b111111111111;
assign Upperletter[208] = 12'b111111111111;
assign Upperletter[209] = 12'b000000000000;
assign Upperletter[210] = 12'b111111111111;
assign Upperletter[211] = 12'b111111111111;
assign Upperletter[212] = 12'b111111111111;
assign Upperletter[213] = 12'b000000000000;
assign Upperletter[214] = 12'b111111111111;
assign Upperletter[215] = 12'b111111111111;
assign Upperletter[216] = 12'b111111111111;
assign Upperletter[217] = 12'b000000000000;
assign Upperletter[218] = 12'b111111111111;
assign Upperletter[219] = 12'b111111111111;
assign Upperletter[220] = 12'b111111111111;
assign Upperletter[221] = 12'b000000000000;
assign Upperletter[222] = 12'b111111111111;
assign Upperletter[223] = 12'b111111111111;
assign Upperletter[224] = 12'b111111111111;
assign Upperletter[225] = 12'b000000000000;
assign Upperletter[226] = 12'b111111111111;
assign Upperletter[227] = 12'b111111111111;
assign Upperletter[228] = 12'b111111111111;
assign Upperletter[229] = 12'b000000000000;
assign Upperletter[230] = 12'b111111111111;
assign Upperletter[231] = 12'b111111111111;
assign Upperletter[232] = 12'b111111111111;
assign Upperletter[233] = 12'b000000000000;
assign Upperletter[234] = 12'b111111111111;
assign Upperletter[235] = 12'b111111111111;
assign Upperletter[236] = 12'b111111111111;
assign Upperletter[237] = 12'b000000000000;
assign Upperletter[238] = 12'b111111111111;
assign Upperletter[239] = 12'b111111111111;
assign Upperletter[240] = 12'b111111111111;
assign Upperletter[241] = 12'b000000000000;
assign Upperletter[242] = 12'b000000000000;
assign Upperletter[243] = 12'b000000000000;
assign Upperletter[244] = 12'b000000000000;
assign Upperletter[245] = 12'b111111111111;
assign Upperletter[246] = 12'b111111111111;
assign Upperletter[247] = 12'b111111111111;
assign Upperletter[248] = 12'b111111111111;
assign Upperletter[249] = 12'b111111111111;
assign Upperletter[250] = 12'b111111111111;
assign Upperletter[251] = 12'b111111111111;
assign Upperletter[252] = 12'b111111111111;
assign Upperletter[253] = 12'b111111111111;
assign Upperletter[254] = 12'b111111111111;
assign Upperletter[255] = 12'b111111111111;
assign Upperletter[256] = 12'b111111111111;
assign Upperletter[257] = 12'b000000000000;
assign Upperletter[258] = 12'b000000000000;
assign Upperletter[259] = 12'b000000000000;
assign Upperletter[260] = 12'b000000000000;
assign Upperletter[261] = 12'b111111111111;
assign Upperletter[262] = 12'b111111111111;
assign Upperletter[263] = 12'b111111111111;
assign Upperletter[264] = 12'b111111111111;
assign Upperletter[265] = 12'b000000000000;
assign Upperletter[266] = 12'b111111111111;
assign Upperletter[267] = 12'b111111111111;
assign Upperletter[268] = 12'b111111111111;
assign Upperletter[269] = 12'b111111111111;
assign Upperletter[270] = 12'b111111111111;
assign Upperletter[271] = 12'b111111111111;
assign Upperletter[272] = 12'b111111111111;
assign Upperletter[273] = 12'b000000000000;
assign Upperletter[274] = 12'b111111111111;
assign Upperletter[275] = 12'b111111111111;
assign Upperletter[276] = 12'b111111111111;
assign Upperletter[277] = 12'b111111111111;
assign Upperletter[278] = 12'b111111111111;
assign Upperletter[279] = 12'b111111111111;
assign Upperletter[280] = 12'b111111111111;
assign Upperletter[281] = 12'b000000000000;
assign Upperletter[282] = 12'b000000000000;
assign Upperletter[283] = 12'b000000000000;
assign Upperletter[284] = 12'b111111111111;
assign Upperletter[285] = 12'b111111111111;
assign Upperletter[286] = 12'b111111111111;
assign Upperletter[287] = 12'b111111111111;
assign Upperletter[288] = 12'b111111111111;
assign Upperletter[289] = 12'b000000000000;
assign Upperletter[290] = 12'b111111111111;
assign Upperletter[291] = 12'b111111111111;
assign Upperletter[292] = 12'b111111111111;
assign Upperletter[293] = 12'b111111111111;
assign Upperletter[294] = 12'b111111111111;
assign Upperletter[295] = 12'b111111111111;
assign Upperletter[296] = 12'b111111111111;
assign Upperletter[297] = 12'b000000000000;
assign Upperletter[298] = 12'b111111111111;
assign Upperletter[299] = 12'b111111111111;
assign Upperletter[300] = 12'b111111111111;
assign Upperletter[301] = 12'b111111111111;
assign Upperletter[302] = 12'b111111111111;
assign Upperletter[303] = 12'b111111111111;
assign Upperletter[304] = 12'b111111111111;
assign Upperletter[305] = 12'b000000000000;
assign Upperletter[306] = 12'b000000000000;
assign Upperletter[307] = 12'b000000000000;
assign Upperletter[308] = 12'b000000000000;
assign Upperletter[309] = 12'b000000000000;
assign Upperletter[310] = 12'b111111111111;
assign Upperletter[311] = 12'b111111111111;
assign Upperletter[312] = 12'b111111111111;
assign Upperletter[313] = 12'b111111111111;
assign Upperletter[314] = 12'b111111111111;
assign Upperletter[315] = 12'b111111111111;
assign Upperletter[316] = 12'b111111111111;
assign Upperletter[317] = 12'b111111111111;
assign Upperletter[318] = 12'b111111111111;
assign Upperletter[319] = 12'b111111111111;
assign Upperletter[320] = 12'b111111111111;
assign Upperletter[321] = 12'b000000000000;
assign Upperletter[322] = 12'b000000000000;
assign Upperletter[323] = 12'b000000000000;
assign Upperletter[324] = 12'b000000000000;
assign Upperletter[325] = 12'b000000000000;
assign Upperletter[326] = 12'b111111111111;
assign Upperletter[327] = 12'b111111111111;
assign Upperletter[328] = 12'b111111111111;
assign Upperletter[329] = 12'b000000000000;
assign Upperletter[330] = 12'b111111111111;
assign Upperletter[331] = 12'b111111111111;
assign Upperletter[332] = 12'b111111111111;
assign Upperletter[333] = 12'b111111111111;
assign Upperletter[334] = 12'b111111111111;
assign Upperletter[335] = 12'b111111111111;
assign Upperletter[336] = 12'b111111111111;
assign Upperletter[337] = 12'b000000000000;
assign Upperletter[338] = 12'b111111111111;
assign Upperletter[339] = 12'b111111111111;
assign Upperletter[340] = 12'b111111111111;
assign Upperletter[341] = 12'b111111111111;
assign Upperletter[342] = 12'b111111111111;
assign Upperletter[343] = 12'b111111111111;
assign Upperletter[344] = 12'b111111111111;
assign Upperletter[345] = 12'b000000000000;
assign Upperletter[346] = 12'b000000000000;
assign Upperletter[347] = 12'b000000000000;
assign Upperletter[348] = 12'b000000000000;
assign Upperletter[349] = 12'b111111111111;
assign Upperletter[350] = 12'b111111111111;
assign Upperletter[351] = 12'b111111111111;
assign Upperletter[352] = 12'b111111111111;
assign Upperletter[353] = 12'b000000000000;
assign Upperletter[354] = 12'b111111111111;
assign Upperletter[355] = 12'b111111111111;
assign Upperletter[356] = 12'b111111111111;
assign Upperletter[357] = 12'b111111111111;
assign Upperletter[358] = 12'b111111111111;
assign Upperletter[359] = 12'b111111111111;
assign Upperletter[360] = 12'b111111111111;
assign Upperletter[361] = 12'b000000000000;
assign Upperletter[362] = 12'b111111111111;
assign Upperletter[363] = 12'b111111111111;
assign Upperletter[364] = 12'b111111111111;
assign Upperletter[365] = 12'b111111111111;
assign Upperletter[366] = 12'b111111111111;
assign Upperletter[367] = 12'b111111111111;
assign Upperletter[368] = 12'b111111111111;
assign Upperletter[369] = 12'b000000000000;
assign Upperletter[370] = 12'b111111111111;
assign Upperletter[371] = 12'b111111111111;
assign Upperletter[372] = 12'b111111111111;
assign Upperletter[373] = 12'b111111111111;
assign Upperletter[374] = 12'b111111111111;
assign Upperletter[375] = 12'b111111111111;
assign Upperletter[376] = 12'b111111111111;
assign Upperletter[377] = 12'b111111111111;
assign Upperletter[378] = 12'b111111111111;
assign Upperletter[379] = 12'b111111111111;
assign Upperletter[380] = 12'b111111111111;
assign Upperletter[381] = 12'b111111111111;
assign Upperletter[382] = 12'b111111111111;
assign Upperletter[383] = 12'b111111111111;
assign Upperletter[384] = 12'b111111111111;
assign Upperletter[385] = 12'b111111111111;
assign Upperletter[386] = 12'b000000000000;
assign Upperletter[387] = 12'b000000000000;
assign Upperletter[388] = 12'b000000000000;
assign Upperletter[389] = 12'b111111111111;
assign Upperletter[390] = 12'b111111111111;
assign Upperletter[391] = 12'b111111111111;
assign Upperletter[392] = 12'b111111111111;
assign Upperletter[393] = 12'b000000000000;
assign Upperletter[394] = 12'b111111111111;
assign Upperletter[395] = 12'b111111111111;
assign Upperletter[396] = 12'b111111111111;
assign Upperletter[397] = 12'b111111111111;
assign Upperletter[398] = 12'b111111111111;
assign Upperletter[399] = 12'b111111111111;
assign Upperletter[400] = 12'b111111111111;
assign Upperletter[401] = 12'b000000000000;
assign Upperletter[402] = 12'b111111111111;
assign Upperletter[403] = 12'b111111111111;
assign Upperletter[404] = 12'b111111111111;
assign Upperletter[405] = 12'b111111111111;
assign Upperletter[406] = 12'b111111111111;
assign Upperletter[407] = 12'b111111111111;
assign Upperletter[408] = 12'b111111111111;
assign Upperletter[409] = 12'b000000000000;
assign Upperletter[410] = 12'b111111111111;
assign Upperletter[411] = 12'b111111111111;
assign Upperletter[412] = 12'b000000000000;
assign Upperletter[413] = 12'b000000000000;
assign Upperletter[414] = 12'b111111111111;
assign Upperletter[415] = 12'b111111111111;
assign Upperletter[416] = 12'b111111111111;
assign Upperletter[417] = 12'b000000000000;
assign Upperletter[418] = 12'b111111111111;
assign Upperletter[419] = 12'b111111111111;
assign Upperletter[420] = 12'b111111111111;
assign Upperletter[421] = 12'b000000000000;
assign Upperletter[422] = 12'b111111111111;
assign Upperletter[423] = 12'b111111111111;
assign Upperletter[424] = 12'b111111111111;
assign Upperletter[425] = 12'b000000000000;
assign Upperletter[426] = 12'b111111111111;
assign Upperletter[427] = 12'b111111111111;
assign Upperletter[428] = 12'b111111111111;
assign Upperletter[429] = 12'b000000000000;
assign Upperletter[430] = 12'b111111111111;
assign Upperletter[431] = 12'b111111111111;
assign Upperletter[432] = 12'b111111111111;
assign Upperletter[433] = 12'b111111111111;
assign Upperletter[434] = 12'b000000000000;
assign Upperletter[435] = 12'b000000000000;
assign Upperletter[436] = 12'b000000000000;
assign Upperletter[437] = 12'b111111111111;
assign Upperletter[438] = 12'b111111111111;
assign Upperletter[439] = 12'b111111111111;
assign Upperletter[440] = 12'b111111111111;
assign Upperletter[441] = 12'b111111111111;
assign Upperletter[442] = 12'b111111111111;
assign Upperletter[443] = 12'b111111111111;
assign Upperletter[444] = 12'b111111111111;
assign Upperletter[445] = 12'b111111111111;
assign Upperletter[446] = 12'b111111111111;
assign Upperletter[447] = 12'b111111111111;
assign Upperletter[448] = 12'b111111111111;
assign Upperletter[449] = 12'b000000000000;
assign Upperletter[450] = 12'b111111111111;
assign Upperletter[451] = 12'b111111111111;
assign Upperletter[452] = 12'b111111111111;
assign Upperletter[453] = 12'b000000000000;
assign Upperletter[454] = 12'b111111111111;
assign Upperletter[455] = 12'b111111111111;
assign Upperletter[456] = 12'b111111111111;
assign Upperletter[457] = 12'b000000000000;
assign Upperletter[458] = 12'b111111111111;
assign Upperletter[459] = 12'b111111111111;
assign Upperletter[460] = 12'b111111111111;
assign Upperletter[461] = 12'b000000000000;
assign Upperletter[462] = 12'b111111111111;
assign Upperletter[463] = 12'b111111111111;
assign Upperletter[464] = 12'b111111111111;
assign Upperletter[465] = 12'b000000000000;
assign Upperletter[466] = 12'b111111111111;
assign Upperletter[467] = 12'b111111111111;
assign Upperletter[468] = 12'b111111111111;
assign Upperletter[469] = 12'b000000000000;
assign Upperletter[470] = 12'b111111111111;
assign Upperletter[471] = 12'b111111111111;
assign Upperletter[472] = 12'b111111111111;
assign Upperletter[473] = 12'b000000000000;
assign Upperletter[474] = 12'b000000000000;
assign Upperletter[475] = 12'b000000000000;
assign Upperletter[476] = 12'b000000000000;
assign Upperletter[477] = 12'b000000000000;
assign Upperletter[478] = 12'b111111111111;
assign Upperletter[479] = 12'b111111111111;
assign Upperletter[480] = 12'b111111111111;
assign Upperletter[481] = 12'b000000000000;
assign Upperletter[482] = 12'b111111111111;
assign Upperletter[483] = 12'b111111111111;
assign Upperletter[484] = 12'b111111111111;
assign Upperletter[485] = 12'b000000000000;
assign Upperletter[486] = 12'b111111111111;
assign Upperletter[487] = 12'b111111111111;
assign Upperletter[488] = 12'b111111111111;
assign Upperletter[489] = 12'b000000000000;
assign Upperletter[490] = 12'b111111111111;
assign Upperletter[491] = 12'b111111111111;
assign Upperletter[492] = 12'b111111111111;
assign Upperletter[493] = 12'b000000000000;
assign Upperletter[494] = 12'b111111111111;
assign Upperletter[495] = 12'b111111111111;
assign Upperletter[496] = 12'b111111111111;
assign Upperletter[497] = 12'b000000000000;
assign Upperletter[498] = 12'b111111111111;
assign Upperletter[499] = 12'b111111111111;
assign Upperletter[500] = 12'b111111111111;
assign Upperletter[501] = 12'b000000000000;
assign Upperletter[502] = 12'b111111111111;
assign Upperletter[503] = 12'b111111111111;
assign Upperletter[504] = 12'b111111111111;
assign Upperletter[505] = 12'b111111111111;
assign Upperletter[506] = 12'b111111111111;
assign Upperletter[507] = 12'b111111111111;
assign Upperletter[508] = 12'b111111111111;
assign Upperletter[509] = 12'b111111111111;
assign Upperletter[510] = 12'b111111111111;
assign Upperletter[511] = 12'b111111111111;
assign Upperletter[512] = 12'b111111111111;
assign Upperletter[513] = 12'b111111111111;
assign Upperletter[514] = 12'b000000000000;
assign Upperletter[515] = 12'b000000000000;
assign Upperletter[516] = 12'b000000000000;
assign Upperletter[517] = 12'b111111111111;
assign Upperletter[518] = 12'b111111111111;
assign Upperletter[519] = 12'b111111111111;
assign Upperletter[520] = 12'b111111111111;
assign Upperletter[521] = 12'b111111111111;
assign Upperletter[522] = 12'b111111111111;
assign Upperletter[523] = 12'b000000000000;
assign Upperletter[524] = 12'b111111111111;
assign Upperletter[525] = 12'b111111111111;
assign Upperletter[526] = 12'b111111111111;
assign Upperletter[527] = 12'b111111111111;
assign Upperletter[528] = 12'b111111111111;
assign Upperletter[529] = 12'b111111111111;
assign Upperletter[530] = 12'b111111111111;
assign Upperletter[531] = 12'b000000000000;
assign Upperletter[532] = 12'b111111111111;
assign Upperletter[533] = 12'b111111111111;
assign Upperletter[534] = 12'b111111111111;
assign Upperletter[535] = 12'b111111111111;
assign Upperletter[536] = 12'b111111111111;
assign Upperletter[537] = 12'b111111111111;
assign Upperletter[538] = 12'b111111111111;
assign Upperletter[539] = 12'b000000000000;
assign Upperletter[540] = 12'b111111111111;
assign Upperletter[541] = 12'b111111111111;
assign Upperletter[542] = 12'b111111111111;
assign Upperletter[543] = 12'b111111111111;
assign Upperletter[544] = 12'b111111111111;
assign Upperletter[545] = 12'b111111111111;
assign Upperletter[546] = 12'b111111111111;
assign Upperletter[547] = 12'b000000000000;
assign Upperletter[548] = 12'b111111111111;
assign Upperletter[549] = 12'b111111111111;
assign Upperletter[550] = 12'b111111111111;
assign Upperletter[551] = 12'b111111111111;
assign Upperletter[552] = 12'b111111111111;
assign Upperletter[553] = 12'b111111111111;
assign Upperletter[554] = 12'b111111111111;
assign Upperletter[555] = 12'b000000000000;
assign Upperletter[556] = 12'b111111111111;
assign Upperletter[557] = 12'b111111111111;
assign Upperletter[558] = 12'b111111111111;
assign Upperletter[559] = 12'b111111111111;
assign Upperletter[560] = 12'b111111111111;
assign Upperletter[561] = 12'b111111111111;
assign Upperletter[562] = 12'b000000000000;
assign Upperletter[563] = 12'b000000000000;
assign Upperletter[564] = 12'b000000000000;
assign Upperletter[565] = 12'b111111111111;
assign Upperletter[566] = 12'b111111111111;
assign Upperletter[567] = 12'b111111111111;
assign Upperletter[568] = 12'b111111111111;
assign Upperletter[569] = 12'b111111111111;
assign Upperletter[570] = 12'b111111111111;
assign Upperletter[571] = 12'b111111111111;
assign Upperletter[572] = 12'b111111111111;
assign Upperletter[573] = 12'b111111111111;
assign Upperletter[574] = 12'b111111111111;
assign Upperletter[575] = 12'b111111111111;
assign Upperletter[576] = 12'b111111111111;
assign Upperletter[577] = 12'b111111111111;
assign Upperletter[578] = 12'b111111111111;
assign Upperletter[579] = 12'b111111111111;
assign Upperletter[580] = 12'b000000000000;
assign Upperletter[581] = 12'b111111111111;
assign Upperletter[582] = 12'b111111111111;
assign Upperletter[583] = 12'b111111111111;
assign Upperletter[584] = 12'b111111111111;
assign Upperletter[585] = 12'b111111111111;
assign Upperletter[586] = 12'b111111111111;
assign Upperletter[587] = 12'b111111111111;
assign Upperletter[588] = 12'b000000000000;
assign Upperletter[589] = 12'b111111111111;
assign Upperletter[590] = 12'b111111111111;
assign Upperletter[591] = 12'b111111111111;
assign Upperletter[592] = 12'b111111111111;
assign Upperletter[593] = 12'b111111111111;
assign Upperletter[594] = 12'b111111111111;
assign Upperletter[595] = 12'b111111111111;
assign Upperletter[596] = 12'b000000000000;
assign Upperletter[597] = 12'b111111111111;
assign Upperletter[598] = 12'b111111111111;
assign Upperletter[599] = 12'b111111111111;
assign Upperletter[600] = 12'b111111111111;
assign Upperletter[601] = 12'b111111111111;
assign Upperletter[602] = 12'b111111111111;
assign Upperletter[603] = 12'b111111111111;
assign Upperletter[604] = 12'b000000000000;
assign Upperletter[605] = 12'b111111111111;
assign Upperletter[606] = 12'b111111111111;
assign Upperletter[607] = 12'b111111111111;
assign Upperletter[608] = 12'b111111111111;
assign Upperletter[609] = 12'b111111111111;
assign Upperletter[610] = 12'b111111111111;
assign Upperletter[611] = 12'b111111111111;
assign Upperletter[612] = 12'b000000000000;
assign Upperletter[613] = 12'b111111111111;
assign Upperletter[614] = 12'b111111111111;
assign Upperletter[615] = 12'b111111111111;
assign Upperletter[616] = 12'b111111111111;
assign Upperletter[617] = 12'b000000000000;
assign Upperletter[618] = 12'b111111111111;
assign Upperletter[619] = 12'b111111111111;
assign Upperletter[620] = 12'b000000000000;
assign Upperletter[621] = 12'b111111111111;
assign Upperletter[622] = 12'b111111111111;
assign Upperletter[623] = 12'b111111111111;
assign Upperletter[624] = 12'b111111111111;
assign Upperletter[625] = 12'b111111111111;
assign Upperletter[626] = 12'b000000000000;
assign Upperletter[627] = 12'b000000000000;
assign Upperletter[628] = 12'b111111111111;
assign Upperletter[629] = 12'b111111111111;
assign Upperletter[630] = 12'b111111111111;
assign Upperletter[631] = 12'b111111111111;
assign Upperletter[632] = 12'b111111111111;
assign Upperletter[633] = 12'b111111111111;
assign Upperletter[634] = 12'b111111111111;
assign Upperletter[635] = 12'b111111111111;
assign Upperletter[636] = 12'b111111111111;
assign Upperletter[637] = 12'b111111111111;
assign Upperletter[638] = 12'b111111111111;
assign Upperletter[639] = 12'b111111111111;
assign Upperletter[640] = 12'b111111111111;
assign Upperletter[641] = 12'b000000000000;
assign Upperletter[642] = 12'b111111111111;
assign Upperletter[643] = 12'b111111111111;
assign Upperletter[644] = 12'b111111111111;
assign Upperletter[645] = 12'b111111111111;
assign Upperletter[646] = 12'b111111111111;
assign Upperletter[647] = 12'b111111111111;
assign Upperletter[648] = 12'b111111111111;
assign Upperletter[649] = 12'b000000000000;
assign Upperletter[650] = 12'b111111111111;
assign Upperletter[651] = 12'b111111111111;
assign Upperletter[652] = 12'b111111111111;
assign Upperletter[653] = 12'b000000000000;
assign Upperletter[654] = 12'b111111111111;
assign Upperletter[655] = 12'b111111111111;
assign Upperletter[656] = 12'b111111111111;
assign Upperletter[657] = 12'b000000000000;
assign Upperletter[658] = 12'b111111111111;
assign Upperletter[659] = 12'b111111111111;
assign Upperletter[660] = 12'b000000000000;
assign Upperletter[661] = 12'b111111111111;
assign Upperletter[662] = 12'b111111111111;
assign Upperletter[663] = 12'b111111111111;
assign Upperletter[664] = 12'b111111111111;
assign Upperletter[665] = 12'b000000000000;
assign Upperletter[666] = 12'b000000000000;
assign Upperletter[667] = 12'b000000000000;
assign Upperletter[668] = 12'b111111111111;
assign Upperletter[669] = 12'b111111111111;
assign Upperletter[670] = 12'b111111111111;
assign Upperletter[671] = 12'b111111111111;
assign Upperletter[672] = 12'b111111111111;
assign Upperletter[673] = 12'b000000000000;
assign Upperletter[674] = 12'b111111111111;
assign Upperletter[675] = 12'b111111111111;
assign Upperletter[676] = 12'b000000000000;
assign Upperletter[677] = 12'b111111111111;
assign Upperletter[678] = 12'b111111111111;
assign Upperletter[679] = 12'b111111111111;
assign Upperletter[680] = 12'b111111111111;
assign Upperletter[681] = 12'b000000000000;
assign Upperletter[682] = 12'b111111111111;
assign Upperletter[683] = 12'b111111111111;
assign Upperletter[684] = 12'b111111111111;
assign Upperletter[685] = 12'b000000000000;
assign Upperletter[686] = 12'b111111111111;
assign Upperletter[687] = 12'b111111111111;
assign Upperletter[688] = 12'b111111111111;
assign Upperletter[689] = 12'b000000000000;
assign Upperletter[690] = 12'b111111111111;
assign Upperletter[691] = 12'b111111111111;
assign Upperletter[692] = 12'b111111111111;
assign Upperletter[693] = 12'b000000000000;
assign Upperletter[694] = 12'b111111111111;
assign Upperletter[695] = 12'b111111111111;
assign Upperletter[696] = 12'b111111111111;
assign Upperletter[697] = 12'b111111111111;
assign Upperletter[698] = 12'b111111111111;
assign Upperletter[699] = 12'b111111111111;
assign Upperletter[700] = 12'b111111111111;
assign Upperletter[701] = 12'b111111111111;
assign Upperletter[702] = 12'b111111111111;
assign Upperletter[703] = 12'b111111111111;
assign Upperletter[704] = 12'b111111111111;
assign Upperletter[705] = 12'b000000000000;
assign Upperletter[706] = 12'b111111111111;
assign Upperletter[707] = 12'b111111111111;
assign Upperletter[708] = 12'b111111111111;
assign Upperletter[709] = 12'b111111111111;
assign Upperletter[710] = 12'b111111111111;
assign Upperletter[711] = 12'b111111111111;
assign Upperletter[712] = 12'b111111111111;
assign Upperletter[713] = 12'b000000000000;
assign Upperletter[714] = 12'b111111111111;
assign Upperletter[715] = 12'b111111111111;
assign Upperletter[716] = 12'b111111111111;
assign Upperletter[717] = 12'b111111111111;
assign Upperletter[718] = 12'b111111111111;
assign Upperletter[719] = 12'b111111111111;
assign Upperletter[720] = 12'b111111111111;
assign Upperletter[721] = 12'b000000000000;
assign Upperletter[722] = 12'b111111111111;
assign Upperletter[723] = 12'b111111111111;
assign Upperletter[724] = 12'b111111111111;
assign Upperletter[725] = 12'b111111111111;
assign Upperletter[726] = 12'b111111111111;
assign Upperletter[727] = 12'b111111111111;
assign Upperletter[728] = 12'b111111111111;
assign Upperletter[729] = 12'b000000000000;
assign Upperletter[730] = 12'b111111111111;
assign Upperletter[731] = 12'b111111111111;
assign Upperletter[732] = 12'b111111111111;
assign Upperletter[733] = 12'b111111111111;
assign Upperletter[734] = 12'b111111111111;
assign Upperletter[735] = 12'b111111111111;
assign Upperletter[736] = 12'b111111111111;
assign Upperletter[737] = 12'b000000000000;
assign Upperletter[738] = 12'b111111111111;
assign Upperletter[739] = 12'b111111111111;
assign Upperletter[740] = 12'b111111111111;
assign Upperletter[741] = 12'b111111111111;
assign Upperletter[742] = 12'b111111111111;
assign Upperletter[743] = 12'b111111111111;
assign Upperletter[744] = 12'b111111111111;
assign Upperletter[745] = 12'b000000000000;
assign Upperletter[746] = 12'b111111111111;
assign Upperletter[747] = 12'b111111111111;
assign Upperletter[748] = 12'b111111111111;
assign Upperletter[749] = 12'b111111111111;
assign Upperletter[750] = 12'b111111111111;
assign Upperletter[751] = 12'b111111111111;
assign Upperletter[752] = 12'b111111111111;
assign Upperletter[753] = 12'b000000000000;
assign Upperletter[754] = 12'b000000000000;
assign Upperletter[755] = 12'b000000000000;
assign Upperletter[756] = 12'b000000000000;
assign Upperletter[757] = 12'b000000000000;
assign Upperletter[758] = 12'b111111111111;
assign Upperletter[759] = 12'b111111111111;
assign Upperletter[760] = 12'b111111111111;
assign Upperletter[761] = 12'b111111111111;
assign Upperletter[762] = 12'b111111111111;
assign Upperletter[763] = 12'b111111111111;
assign Upperletter[764] = 12'b111111111111;
assign Upperletter[765] = 12'b111111111111;
assign Upperletter[766] = 12'b111111111111;
assign Upperletter[767] = 12'b111111111111;
assign Upperletter[768] = 12'b111111111111;
assign Upperletter[769] = 12'b000000000000;
assign Upperletter[770] = 12'b111111111111;
assign Upperletter[771] = 12'b111111111111;
assign Upperletter[772] = 12'b111111111111;
assign Upperletter[773] = 12'b000000000000;
assign Upperletter[774] = 12'b111111111111;
assign Upperletter[775] = 12'b111111111111;
assign Upperletter[776] = 12'b111111111111;
assign Upperletter[777] = 12'b000000000000;
assign Upperletter[778] = 12'b000000000000;
assign Upperletter[779] = 12'b111111111111;
assign Upperletter[780] = 12'b000000000000;
assign Upperletter[781] = 12'b000000000000;
assign Upperletter[782] = 12'b111111111111;
assign Upperletter[783] = 12'b111111111111;
assign Upperletter[784] = 12'b111111111111;
assign Upperletter[785] = 12'b000000000000;
assign Upperletter[786] = 12'b111111111111;
assign Upperletter[787] = 12'b000000000000;
assign Upperletter[788] = 12'b111111111111;
assign Upperletter[789] = 12'b000000000000;
assign Upperletter[790] = 12'b111111111111;
assign Upperletter[791] = 12'b111111111111;
assign Upperletter[792] = 12'b111111111111;
assign Upperletter[793] = 12'b000000000000;
assign Upperletter[794] = 12'b111111111111;
assign Upperletter[795] = 12'b111111111111;
assign Upperletter[796] = 12'b111111111111;
assign Upperletter[797] = 12'b000000000000;
assign Upperletter[798] = 12'b111111111111;
assign Upperletter[799] = 12'b111111111111;
assign Upperletter[800] = 12'b111111111111;
assign Upperletter[801] = 12'b000000000000;
assign Upperletter[802] = 12'b111111111111;
assign Upperletter[803] = 12'b111111111111;
assign Upperletter[804] = 12'b111111111111;
assign Upperletter[805] = 12'b000000000000;
assign Upperletter[806] = 12'b111111111111;
assign Upperletter[807] = 12'b111111111111;
assign Upperletter[808] = 12'b111111111111;
assign Upperletter[809] = 12'b000000000000;
assign Upperletter[810] = 12'b111111111111;
assign Upperletter[811] = 12'b111111111111;
assign Upperletter[812] = 12'b111111111111;
assign Upperletter[813] = 12'b000000000000;
assign Upperletter[814] = 12'b111111111111;
assign Upperletter[815] = 12'b111111111111;
assign Upperletter[816] = 12'b111111111111;
assign Upperletter[817] = 12'b000000000000;
assign Upperletter[818] = 12'b111111111111;
assign Upperletter[819] = 12'b111111111111;
assign Upperletter[820] = 12'b111111111111;
assign Upperletter[821] = 12'b000000000000;
assign Upperletter[822] = 12'b111111111111;
assign Upperletter[823] = 12'b111111111111;
assign Upperletter[824] = 12'b111111111111;
assign Upperletter[825] = 12'b111111111111;
assign Upperletter[826] = 12'b111111111111;
assign Upperletter[827] = 12'b111111111111;
assign Upperletter[828] = 12'b111111111111;
assign Upperletter[829] = 12'b111111111111;
assign Upperletter[830] = 12'b111111111111;
assign Upperletter[831] = 12'b111111111111;
assign Upperletter[832] = 12'b111111111111;
assign Upperletter[833] = 12'b000000000000;
assign Upperletter[834] = 12'b111111111111;
assign Upperletter[835] = 12'b111111111111;
assign Upperletter[836] = 12'b111111111111;
assign Upperletter[837] = 12'b000000000000;
assign Upperletter[838] = 12'b111111111111;
assign Upperletter[839] = 12'b111111111111;
assign Upperletter[840] = 12'b111111111111;
assign Upperletter[841] = 12'b000000000000;
assign Upperletter[842] = 12'b000000000000;
assign Upperletter[843] = 12'b111111111111;
assign Upperletter[844] = 12'b111111111111;
assign Upperletter[845] = 12'b000000000000;
assign Upperletter[846] = 12'b111111111111;
assign Upperletter[847] = 12'b111111111111;
assign Upperletter[848] = 12'b111111111111;
assign Upperletter[849] = 12'b000000000000;
assign Upperletter[850] = 12'b111111111111;
assign Upperletter[851] = 12'b000000000000;
assign Upperletter[852] = 12'b111111111111;
assign Upperletter[853] = 12'b000000000000;
assign Upperletter[854] = 12'b111111111111;
assign Upperletter[855] = 12'b111111111111;
assign Upperletter[856] = 12'b111111111111;
assign Upperletter[857] = 12'b000000000000;
assign Upperletter[858] = 12'b111111111111;
assign Upperletter[859] = 12'b111111111111;
assign Upperletter[860] = 12'b000000000000;
assign Upperletter[861] = 12'b000000000000;
assign Upperletter[862] = 12'b111111111111;
assign Upperletter[863] = 12'b111111111111;
assign Upperletter[864] = 12'b111111111111;
assign Upperletter[865] = 12'b000000000000;
assign Upperletter[866] = 12'b111111111111;
assign Upperletter[867] = 12'b111111111111;
assign Upperletter[868] = 12'b111111111111;
assign Upperletter[869] = 12'b000000000000;
assign Upperletter[870] = 12'b111111111111;
assign Upperletter[871] = 12'b111111111111;
assign Upperletter[872] = 12'b111111111111;
assign Upperletter[873] = 12'b000000000000;
assign Upperletter[874] = 12'b111111111111;
assign Upperletter[875] = 12'b111111111111;
assign Upperletter[876] = 12'b111111111111;
assign Upperletter[877] = 12'b000000000000;
assign Upperletter[878] = 12'b111111111111;
assign Upperletter[879] = 12'b111111111111;
assign Upperletter[880] = 12'b111111111111;
assign Upperletter[881] = 12'b000000000000;
assign Upperletter[882] = 12'b111111111111;
assign Upperletter[883] = 12'b111111111111;
assign Upperletter[884] = 12'b111111111111;
assign Upperletter[885] = 12'b000000000000;
assign Upperletter[886] = 12'b111111111111;
assign Upperletter[887] = 12'b111111111111;
assign Upperletter[888] = 12'b111111111111;
assign Upperletter[889] = 12'b111111111111;
assign Upperletter[890] = 12'b111111111111;
assign Upperletter[891] = 12'b111111111111;
assign Upperletter[892] = 12'b111111111111;
assign Upperletter[893] = 12'b111111111111;
assign Upperletter[894] = 12'b111111111111;
assign Upperletter[895] = 12'b111111111111;
assign Upperletter[896] = 12'b111111111111;
assign Upperletter[897] = 12'b111111111111;
assign Upperletter[898] = 12'b000000000000;
assign Upperletter[899] = 12'b000000000000;
assign Upperletter[900] = 12'b000000000000;
assign Upperletter[901] = 12'b111111111111;
assign Upperletter[902] = 12'b111111111111;
assign Upperletter[903] = 12'b111111111111;
assign Upperletter[904] = 12'b111111111111;
assign Upperletter[905] = 12'b000000000000;
assign Upperletter[906] = 12'b111111111111;
assign Upperletter[907] = 12'b111111111111;
assign Upperletter[908] = 12'b111111111111;
assign Upperletter[909] = 12'b000000000000;
assign Upperletter[910] = 12'b111111111111;
assign Upperletter[911] = 12'b111111111111;
assign Upperletter[912] = 12'b111111111111;
assign Upperletter[913] = 12'b000000000000;
assign Upperletter[914] = 12'b111111111111;
assign Upperletter[915] = 12'b111111111111;
assign Upperletter[916] = 12'b111111111111;
assign Upperletter[917] = 12'b000000000000;
assign Upperletter[918] = 12'b111111111111;
assign Upperletter[919] = 12'b111111111111;
assign Upperletter[920] = 12'b111111111111;
assign Upperletter[921] = 12'b000000000000;
assign Upperletter[922] = 12'b111111111111;
assign Upperletter[923] = 12'b111111111111;
assign Upperletter[924] = 12'b111111111111;
assign Upperletter[925] = 12'b000000000000;
assign Upperletter[926] = 12'b111111111111;
assign Upperletter[927] = 12'b111111111111;
assign Upperletter[928] = 12'b111111111111;
assign Upperletter[929] = 12'b000000000000;
assign Upperletter[930] = 12'b111111111111;
assign Upperletter[931] = 12'b111111111111;
assign Upperletter[932] = 12'b111111111111;
assign Upperletter[933] = 12'b000000000000;
assign Upperletter[934] = 12'b111111111111;
assign Upperletter[935] = 12'b111111111111;
assign Upperletter[936] = 12'b111111111111;
assign Upperletter[937] = 12'b000000000000;
assign Upperletter[938] = 12'b111111111111;
assign Upperletter[939] = 12'b111111111111;
assign Upperletter[940] = 12'b111111111111;
assign Upperletter[941] = 12'b000000000000;
assign Upperletter[942] = 12'b111111111111;
assign Upperletter[943] = 12'b111111111111;
assign Upperletter[944] = 12'b111111111111;
assign Upperletter[945] = 12'b111111111111;
assign Upperletter[946] = 12'b000000000000;
assign Upperletter[947] = 12'b000000000000;
assign Upperletter[948] = 12'b000000000000;
assign Upperletter[949] = 12'b111111111111;
assign Upperletter[950] = 12'b111111111111;
assign Upperletter[951] = 12'b111111111111;
assign Upperletter[952] = 12'b111111111111;
assign Upperletter[953] = 12'b111111111111;
assign Upperletter[954] = 12'b111111111111;
assign Upperletter[955] = 12'b111111111111;
assign Upperletter[956] = 12'b111111111111;
assign Upperletter[957] = 12'b111111111111;
assign Upperletter[958] = 12'b111111111111;
assign Upperletter[959] = 12'b111111111111;
assign Upperletter[960] = 12'b111111111111;
assign Upperletter[961] = 12'b000000000000;
assign Upperletter[962] = 12'b000000000000;
assign Upperletter[963] = 12'b000000000000;
assign Upperletter[964] = 12'b000000000000;
assign Upperletter[965] = 12'b111111111111;
assign Upperletter[966] = 12'b111111111111;
assign Upperletter[967] = 12'b111111111111;
assign Upperletter[968] = 12'b111111111111;
assign Upperletter[969] = 12'b000000000000;
assign Upperletter[970] = 12'b111111111111;
assign Upperletter[971] = 12'b111111111111;
assign Upperletter[972] = 12'b111111111111;
assign Upperletter[973] = 12'b000000000000;
assign Upperletter[974] = 12'b111111111111;
assign Upperletter[975] = 12'b111111111111;
assign Upperletter[976] = 12'b111111111111;
assign Upperletter[977] = 12'b000000000000;
assign Upperletter[978] = 12'b111111111111;
assign Upperletter[979] = 12'b111111111111;
assign Upperletter[980] = 12'b111111111111;
assign Upperletter[981] = 12'b000000000000;
assign Upperletter[982] = 12'b111111111111;
assign Upperletter[983] = 12'b111111111111;
assign Upperletter[984] = 12'b111111111111;
assign Upperletter[985] = 12'b000000000000;
assign Upperletter[986] = 12'b000000000000;
assign Upperletter[987] = 12'b000000000000;
assign Upperletter[988] = 12'b000000000000;
assign Upperletter[989] = 12'b111111111111;
assign Upperletter[990] = 12'b111111111111;
assign Upperletter[991] = 12'b111111111111;
assign Upperletter[992] = 12'b111111111111;
assign Upperletter[993] = 12'b000000000000;
assign Upperletter[994] = 12'b111111111111;
assign Upperletter[995] = 12'b111111111111;
assign Upperletter[996] = 12'b111111111111;
assign Upperletter[997] = 12'b111111111111;
assign Upperletter[998] = 12'b111111111111;
assign Upperletter[999] = 12'b111111111111;
assign Upperletter[1000] = 12'b111111111111;
assign Upperletter[1001] = 12'b000000000000;
assign Upperletter[1002] = 12'b111111111111;
assign Upperletter[1003] = 12'b111111111111;
assign Upperletter[1004] = 12'b111111111111;
assign Upperletter[1005] = 12'b111111111111;
assign Upperletter[1006] = 12'b111111111111;
assign Upperletter[1007] = 12'b111111111111;
assign Upperletter[1008] = 12'b111111111111;
assign Upperletter[1009] = 12'b000000000000;
assign Upperletter[1010] = 12'b111111111111;
assign Upperletter[1011] = 12'b111111111111;
assign Upperletter[1012] = 12'b111111111111;
assign Upperletter[1013] = 12'b111111111111;
assign Upperletter[1014] = 12'b111111111111;
assign Upperletter[1015] = 12'b111111111111;
assign Upperletter[1016] = 12'b111111111111;
assign Upperletter[1017] = 12'b111111111111;
assign Upperletter[1018] = 12'b111111111111;
assign Upperletter[1019] = 12'b111111111111;
assign Upperletter[1020] = 12'b111111111111;
assign Upperletter[1021] = 12'b111111111111;
assign Upperletter[1022] = 12'b111111111111;
assign Upperletter[1023] = 12'b111111111111;
assign Upperletter[1024] = 12'b111111111111;
assign Upperletter[1025] = 12'b111111111111;
assign Upperletter[1026] = 12'b000000000000;
assign Upperletter[1027] = 12'b000000000000;
assign Upperletter[1028] = 12'b000000000000;
assign Upperletter[1029] = 12'b111111111111;
assign Upperletter[1030] = 12'b111111111111;
assign Upperletter[1031] = 12'b111111111111;
assign Upperletter[1032] = 12'b111111111111;
assign Upperletter[1033] = 12'b000000000000;
assign Upperletter[1034] = 12'b111111111111;
assign Upperletter[1035] = 12'b111111111111;
assign Upperletter[1036] = 12'b111111111111;
assign Upperletter[1037] = 12'b000000000000;
assign Upperletter[1038] = 12'b111111111111;
assign Upperletter[1039] = 12'b111111111111;
assign Upperletter[1040] = 12'b111111111111;
assign Upperletter[1041] = 12'b000000000000;
assign Upperletter[1042] = 12'b111111111111;
assign Upperletter[1043] = 12'b111111111111;
assign Upperletter[1044] = 12'b111111111111;
assign Upperletter[1045] = 12'b000000000000;
assign Upperletter[1046] = 12'b111111111111;
assign Upperletter[1047] = 12'b111111111111;
assign Upperletter[1048] = 12'b111111111111;
assign Upperletter[1049] = 12'b000000000000;
assign Upperletter[1050] = 12'b111111111111;
assign Upperletter[1051] = 12'b111111111111;
assign Upperletter[1052] = 12'b111111111111;
assign Upperletter[1053] = 12'b000000000000;
assign Upperletter[1054] = 12'b111111111111;
assign Upperletter[1055] = 12'b111111111111;
assign Upperletter[1056] = 12'b111111111111;
assign Upperletter[1057] = 12'b000000000000;
assign Upperletter[1058] = 12'b111111111111;
assign Upperletter[1059] = 12'b111111111111;
assign Upperletter[1060] = 12'b111111111111;
assign Upperletter[1061] = 12'b000000000000;
assign Upperletter[1062] = 12'b111111111111;
assign Upperletter[1063] = 12'b111111111111;
assign Upperletter[1064] = 12'b111111111111;
assign Upperletter[1065] = 12'b000000000000;
assign Upperletter[1066] = 12'b111111111111;
assign Upperletter[1067] = 12'b111111111111;
assign Upperletter[1068] = 12'b000000000000;
assign Upperletter[1069] = 12'b111111111111;
assign Upperletter[1070] = 12'b111111111111;
assign Upperletter[1071] = 12'b111111111111;
assign Upperletter[1072] = 12'b111111111111;
assign Upperletter[1073] = 12'b111111111111;
assign Upperletter[1074] = 12'b000000000000;
assign Upperletter[1075] = 12'b000000000000;
assign Upperletter[1076] = 12'b111111111111;
assign Upperletter[1077] = 12'b000000000000;
assign Upperletter[1078] = 12'b111111111111;
assign Upperletter[1079] = 12'b111111111111;
assign Upperletter[1080] = 12'b111111111111;
assign Upperletter[1081] = 12'b111111111111;
assign Upperletter[1082] = 12'b111111111111;
assign Upperletter[1083] = 12'b111111111111;
assign Upperletter[1084] = 12'b111111111111;
assign Upperletter[1085] = 12'b111111111111;
assign Upperletter[1086] = 12'b111111111111;
assign Upperletter[1087] = 12'b111111111111;
assign Upperletter[1088] = 12'b111111111111;
assign Upperletter[1089] = 12'b000000000000;
assign Upperletter[1090] = 12'b000000000000;
assign Upperletter[1091] = 12'b000000000000;
assign Upperletter[1092] = 12'b000000000000;
assign Upperletter[1093] = 12'b111111111111;
assign Upperletter[1094] = 12'b111111111111;
assign Upperletter[1095] = 12'b111111111111;
assign Upperletter[1096] = 12'b111111111111;
assign Upperletter[1097] = 12'b000000000000;
assign Upperletter[1098] = 12'b111111111111;
assign Upperletter[1099] = 12'b111111111111;
assign Upperletter[1100] = 12'b111111111111;
assign Upperletter[1101] = 12'b000000000000;
assign Upperletter[1102] = 12'b111111111111;
assign Upperletter[1103] = 12'b111111111111;
assign Upperletter[1104] = 12'b111111111111;
assign Upperletter[1105] = 12'b000000000000;
assign Upperletter[1106] = 12'b111111111111;
assign Upperletter[1107] = 12'b111111111111;
assign Upperletter[1108] = 12'b111111111111;
assign Upperletter[1109] = 12'b000000000000;
assign Upperletter[1110] = 12'b111111111111;
assign Upperletter[1111] = 12'b111111111111;
assign Upperletter[1112] = 12'b111111111111;
assign Upperletter[1113] = 12'b000000000000;
assign Upperletter[1114] = 12'b000000000000;
assign Upperletter[1115] = 12'b000000000000;
assign Upperletter[1116] = 12'b000000000000;
assign Upperletter[1117] = 12'b111111111111;
assign Upperletter[1118] = 12'b111111111111;
assign Upperletter[1119] = 12'b111111111111;
assign Upperletter[1120] = 12'b111111111111;
assign Upperletter[1121] = 12'b000000000000;
assign Upperletter[1122] = 12'b111111111111;
assign Upperletter[1123] = 12'b000000000000;
assign Upperletter[1124] = 12'b111111111111;
assign Upperletter[1125] = 12'b111111111111;
assign Upperletter[1126] = 12'b111111111111;
assign Upperletter[1127] = 12'b111111111111;
assign Upperletter[1128] = 12'b111111111111;
assign Upperletter[1129] = 12'b000000000000;
assign Upperletter[1130] = 12'b111111111111;
assign Upperletter[1131] = 12'b111111111111;
assign Upperletter[1132] = 12'b000000000000;
assign Upperletter[1133] = 12'b111111111111;
assign Upperletter[1134] = 12'b111111111111;
assign Upperletter[1135] = 12'b111111111111;
assign Upperletter[1136] = 12'b111111111111;
assign Upperletter[1137] = 12'b000000000000;
assign Upperletter[1138] = 12'b111111111111;
assign Upperletter[1139] = 12'b111111111111;
assign Upperletter[1140] = 12'b111111111111;
assign Upperletter[1141] = 12'b000000000000;
assign Upperletter[1142] = 12'b111111111111;
assign Upperletter[1143] = 12'b111111111111;
assign Upperletter[1144] = 12'b111111111111;
assign Upperletter[1145] = 12'b111111111111;
assign Upperletter[1146] = 12'b111111111111;
assign Upperletter[1147] = 12'b111111111111;
assign Upperletter[1148] = 12'b111111111111;
assign Upperletter[1149] = 12'b111111111111;
assign Upperletter[1150] = 12'b111111111111;
assign Upperletter[1151] = 12'b111111111111;
assign Upperletter[1152] = 12'b111111111111;
assign Upperletter[1153] = 12'b111111111111;
assign Upperletter[1154] = 12'b000000000000;
assign Upperletter[1155] = 12'b000000000000;
assign Upperletter[1156] = 12'b000000000000;
assign Upperletter[1157] = 12'b000000000000;
assign Upperletter[1158] = 12'b111111111111;
assign Upperletter[1159] = 12'b111111111111;
assign Upperletter[1160] = 12'b111111111111;
assign Upperletter[1161] = 12'b000000000000;
assign Upperletter[1162] = 12'b111111111111;
assign Upperletter[1163] = 12'b111111111111;
assign Upperletter[1164] = 12'b111111111111;
assign Upperletter[1165] = 12'b111111111111;
assign Upperletter[1166] = 12'b111111111111;
assign Upperletter[1167] = 12'b111111111111;
assign Upperletter[1168] = 12'b111111111111;
assign Upperletter[1169] = 12'b000000000000;
assign Upperletter[1170] = 12'b111111111111;
assign Upperletter[1171] = 12'b111111111111;
assign Upperletter[1172] = 12'b111111111111;
assign Upperletter[1173] = 12'b111111111111;
assign Upperletter[1174] = 12'b111111111111;
assign Upperletter[1175] = 12'b111111111111;
assign Upperletter[1176] = 12'b111111111111;
assign Upperletter[1177] = 12'b111111111111;
assign Upperletter[1178] = 12'b000000000000;
assign Upperletter[1179] = 12'b000000000000;
assign Upperletter[1180] = 12'b000000000000;
assign Upperletter[1181] = 12'b111111111111;
assign Upperletter[1182] = 12'b111111111111;
assign Upperletter[1183] = 12'b111111111111;
assign Upperletter[1184] = 12'b111111111111;
assign Upperletter[1185] = 12'b111111111111;
assign Upperletter[1186] = 12'b111111111111;
assign Upperletter[1187] = 12'b111111111111;
assign Upperletter[1188] = 12'b111111111111;
assign Upperletter[1189] = 12'b000000000000;
assign Upperletter[1190] = 12'b111111111111;
assign Upperletter[1191] = 12'b111111111111;
assign Upperletter[1192] = 12'b111111111111;
assign Upperletter[1193] = 12'b111111111111;
assign Upperletter[1194] = 12'b111111111111;
assign Upperletter[1195] = 12'b111111111111;
assign Upperletter[1196] = 12'b111111111111;
assign Upperletter[1197] = 12'b000000000000;
assign Upperletter[1198] = 12'b111111111111;
assign Upperletter[1199] = 12'b111111111111;
assign Upperletter[1200] = 12'b111111111111;
assign Upperletter[1201] = 12'b000000000000;
assign Upperletter[1202] = 12'b000000000000;
assign Upperletter[1203] = 12'b000000000000;
assign Upperletter[1204] = 12'b000000000000;
assign Upperletter[1205] = 12'b111111111111;
assign Upperletter[1206] = 12'b111111111111;
assign Upperletter[1207] = 12'b111111111111;
assign Upperletter[1208] = 12'b111111111111;
assign Upperletter[1209] = 12'b111111111111;
assign Upperletter[1210] = 12'b111111111111;
assign Upperletter[1211] = 12'b111111111111;
assign Upperletter[1212] = 12'b111111111111;
assign Upperletter[1213] = 12'b111111111111;
assign Upperletter[1214] = 12'b111111111111;
assign Upperletter[1215] = 12'b111111111111;
assign Upperletter[1216] = 12'b111111111111;
assign Upperletter[1217] = 12'b000000000000;
assign Upperletter[1218] = 12'b000000000000;
assign Upperletter[1219] = 12'b000000000000;
assign Upperletter[1220] = 12'b000000000000;
assign Upperletter[1221] = 12'b000000000000;
assign Upperletter[1222] = 12'b111111111111;
assign Upperletter[1223] = 12'b111111111111;
assign Upperletter[1224] = 12'b111111111111;
assign Upperletter[1225] = 12'b111111111111;
assign Upperletter[1226] = 12'b111111111111;
assign Upperletter[1227] = 12'b000000000000;
assign Upperletter[1228] = 12'b111111111111;
assign Upperletter[1229] = 12'b111111111111;
assign Upperletter[1230] = 12'b111111111111;
assign Upperletter[1231] = 12'b111111111111;
assign Upperletter[1232] = 12'b111111111111;
assign Upperletter[1233] = 12'b111111111111;
assign Upperletter[1234] = 12'b111111111111;
assign Upperletter[1235] = 12'b000000000000;
assign Upperletter[1236] = 12'b111111111111;
assign Upperletter[1237] = 12'b111111111111;
assign Upperletter[1238] = 12'b111111111111;
assign Upperletter[1239] = 12'b111111111111;
assign Upperletter[1240] = 12'b111111111111;
assign Upperletter[1241] = 12'b111111111111;
assign Upperletter[1242] = 12'b111111111111;
assign Upperletter[1243] = 12'b000000000000;
assign Upperletter[1244] = 12'b111111111111;
assign Upperletter[1245] = 12'b111111111111;
assign Upperletter[1246] = 12'b111111111111;
assign Upperletter[1247] = 12'b111111111111;
assign Upperletter[1248] = 12'b111111111111;
assign Upperletter[1249] = 12'b111111111111;
assign Upperletter[1250] = 12'b111111111111;
assign Upperletter[1251] = 12'b000000000000;
assign Upperletter[1252] = 12'b111111111111;
assign Upperletter[1253] = 12'b111111111111;
assign Upperletter[1254] = 12'b111111111111;
assign Upperletter[1255] = 12'b111111111111;
assign Upperletter[1256] = 12'b111111111111;
assign Upperletter[1257] = 12'b111111111111;
assign Upperletter[1258] = 12'b111111111111;
assign Upperletter[1259] = 12'b000000000000;
assign Upperletter[1260] = 12'b111111111111;
assign Upperletter[1261] = 12'b111111111111;
assign Upperletter[1262] = 12'b111111111111;
assign Upperletter[1263] = 12'b111111111111;
assign Upperletter[1264] = 12'b111111111111;
assign Upperletter[1265] = 12'b111111111111;
assign Upperletter[1266] = 12'b111111111111;
assign Upperletter[1267] = 12'b000000000000;
assign Upperletter[1268] = 12'b111111111111;
assign Upperletter[1269] = 12'b111111111111;
assign Upperletter[1270] = 12'b111111111111;
assign Upperletter[1271] = 12'b111111111111;
assign Upperletter[1272] = 12'b111111111111;
assign Upperletter[1273] = 12'b111111111111;
assign Upperletter[1274] = 12'b111111111111;
assign Upperletter[1275] = 12'b111111111111;
assign Upperletter[1276] = 12'b111111111111;
assign Upperletter[1277] = 12'b111111111111;
assign Upperletter[1278] = 12'b111111111111;
assign Upperletter[1279] = 12'b111111111111;
assign Upperletter[1280] = 12'b111111111111;
assign Upperletter[1281] = 12'b000000000000;
assign Upperletter[1282] = 12'b111111111111;
assign Upperletter[1283] = 12'b111111111111;
assign Upperletter[1284] = 12'b111111111111;
assign Upperletter[1285] = 12'b000000000000;
assign Upperletter[1286] = 12'b111111111111;
assign Upperletter[1287] = 12'b111111111111;
assign Upperletter[1288] = 12'b111111111111;
assign Upperletter[1289] = 12'b000000000000;
assign Upperletter[1290] = 12'b111111111111;
assign Upperletter[1291] = 12'b111111111111;
assign Upperletter[1292] = 12'b111111111111;
assign Upperletter[1293] = 12'b000000000000;
assign Upperletter[1294] = 12'b111111111111;
assign Upperletter[1295] = 12'b111111111111;
assign Upperletter[1296] = 12'b111111111111;
assign Upperletter[1297] = 12'b000000000000;
assign Upperletter[1298] = 12'b111111111111;
assign Upperletter[1299] = 12'b111111111111;
assign Upperletter[1300] = 12'b111111111111;
assign Upperletter[1301] = 12'b000000000000;
assign Upperletter[1302] = 12'b111111111111;
assign Upperletter[1303] = 12'b111111111111;
assign Upperletter[1304] = 12'b111111111111;
assign Upperletter[1305] = 12'b000000000000;
assign Upperletter[1306] = 12'b111111111111;
assign Upperletter[1307] = 12'b111111111111;
assign Upperletter[1308] = 12'b111111111111;
assign Upperletter[1309] = 12'b000000000000;
assign Upperletter[1310] = 12'b111111111111;
assign Upperletter[1311] = 12'b111111111111;
assign Upperletter[1312] = 12'b111111111111;
assign Upperletter[1313] = 12'b000000000000;
assign Upperletter[1314] = 12'b111111111111;
assign Upperletter[1315] = 12'b111111111111;
assign Upperletter[1316] = 12'b111111111111;
assign Upperletter[1317] = 12'b000000000000;
assign Upperletter[1318] = 12'b111111111111;
assign Upperletter[1319] = 12'b111111111111;
assign Upperletter[1320] = 12'b111111111111;
assign Upperletter[1321] = 12'b000000000000;
assign Upperletter[1322] = 12'b111111111111;
assign Upperletter[1323] = 12'b111111111111;
assign Upperletter[1324] = 12'b111111111111;
assign Upperletter[1325] = 12'b000000000000;
assign Upperletter[1326] = 12'b111111111111;
assign Upperletter[1327] = 12'b111111111111;
assign Upperletter[1328] = 12'b111111111111;
assign Upperletter[1329] = 12'b111111111111;
assign Upperletter[1330] = 12'b000000000000;
assign Upperletter[1331] = 12'b000000000000;
assign Upperletter[1332] = 12'b000000000000;
assign Upperletter[1333] = 12'b111111111111;
assign Upperletter[1334] = 12'b111111111111;
assign Upperletter[1335] = 12'b111111111111;
assign Upperletter[1336] = 12'b111111111111;
assign Upperletter[1337] = 12'b111111111111;
assign Upperletter[1338] = 12'b111111111111;
assign Upperletter[1339] = 12'b111111111111;
assign Upperletter[1340] = 12'b111111111111;
assign Upperletter[1341] = 12'b111111111111;
assign Upperletter[1342] = 12'b111111111111;
assign Upperletter[1343] = 12'b111111111111;
assign Upperletter[1344] = 12'b111111111111;
assign Upperletter[1345] = 12'b000000000000;
assign Upperletter[1346] = 12'b111111111111;
assign Upperletter[1347] = 12'b111111111111;
assign Upperletter[1348] = 12'b111111111111;
assign Upperletter[1349] = 12'b000000000000;
assign Upperletter[1350] = 12'b111111111111;
assign Upperletter[1351] = 12'b111111111111;
assign Upperletter[1352] = 12'b111111111111;
assign Upperletter[1353] = 12'b000000000000;
assign Upperletter[1354] = 12'b111111111111;
assign Upperletter[1355] = 12'b111111111111;
assign Upperletter[1356] = 12'b111111111111;
assign Upperletter[1357] = 12'b000000000000;
assign Upperletter[1358] = 12'b111111111111;
assign Upperletter[1359] = 12'b111111111111;
assign Upperletter[1360] = 12'b111111111111;
assign Upperletter[1361] = 12'b000000000000;
assign Upperletter[1362] = 12'b111111111111;
assign Upperletter[1363] = 12'b111111111111;
assign Upperletter[1364] = 12'b111111111111;
assign Upperletter[1365] = 12'b000000000000;
assign Upperletter[1366] = 12'b111111111111;
assign Upperletter[1367] = 12'b111111111111;
assign Upperletter[1368] = 12'b111111111111;
assign Upperletter[1369] = 12'b000000000000;
assign Upperletter[1370] = 12'b111111111111;
assign Upperletter[1371] = 12'b111111111111;
assign Upperletter[1372] = 12'b111111111111;
assign Upperletter[1373] = 12'b000000000000;
assign Upperletter[1374] = 12'b111111111111;
assign Upperletter[1375] = 12'b111111111111;
assign Upperletter[1376] = 12'b111111111111;
assign Upperletter[1377] = 12'b000000000000;
assign Upperletter[1378] = 12'b111111111111;
assign Upperletter[1379] = 12'b111111111111;
assign Upperletter[1380] = 12'b111111111111;
assign Upperletter[1381] = 12'b000000000000;
assign Upperletter[1382] = 12'b111111111111;
assign Upperletter[1383] = 12'b111111111111;
assign Upperletter[1384] = 12'b111111111111;
assign Upperletter[1385] = 12'b111111111111;
assign Upperletter[1386] = 12'b000000000000;
assign Upperletter[1387] = 12'b111111111111;
assign Upperletter[1388] = 12'b000000000000;
assign Upperletter[1389] = 12'b111111111111;
assign Upperletter[1390] = 12'b111111111111;
assign Upperletter[1391] = 12'b111111111111;
assign Upperletter[1392] = 12'b111111111111;
assign Upperletter[1393] = 12'b111111111111;
assign Upperletter[1394] = 12'b111111111111;
assign Upperletter[1395] = 12'b000000000000;
assign Upperletter[1396] = 12'b111111111111;
assign Upperletter[1397] = 12'b111111111111;
assign Upperletter[1398] = 12'b111111111111;
assign Upperletter[1399] = 12'b111111111111;
assign Upperletter[1400] = 12'b111111111111;
assign Upperletter[1401] = 12'b111111111111;
assign Upperletter[1402] = 12'b111111111111;
assign Upperletter[1403] = 12'b111111111111;
assign Upperletter[1404] = 12'b111111111111;
assign Upperletter[1405] = 12'b111111111111;
assign Upperletter[1406] = 12'b111111111111;
assign Upperletter[1407] = 12'b111111111111;
assign Upperletter[1408] = 12'b111111111111;
assign Upperletter[1409] = 12'b000000000000;
assign Upperletter[1410] = 12'b111111111111;
assign Upperletter[1411] = 12'b111111111111;
assign Upperletter[1412] = 12'b111111111111;
assign Upperletter[1413] = 12'b000000000000;
assign Upperletter[1414] = 12'b111111111111;
assign Upperletter[1415] = 12'b111111111111;
assign Upperletter[1416] = 12'b111111111111;
assign Upperletter[1417] = 12'b000000000000;
assign Upperletter[1418] = 12'b111111111111;
assign Upperletter[1419] = 12'b111111111111;
assign Upperletter[1420] = 12'b111111111111;
assign Upperletter[1421] = 12'b000000000000;
assign Upperletter[1422] = 12'b111111111111;
assign Upperletter[1423] = 12'b111111111111;
assign Upperletter[1424] = 12'b111111111111;
assign Upperletter[1425] = 12'b000000000000;
assign Upperletter[1426] = 12'b111111111111;
assign Upperletter[1427] = 12'b111111111111;
assign Upperletter[1428] = 12'b111111111111;
assign Upperletter[1429] = 12'b000000000000;
assign Upperletter[1430] = 12'b111111111111;
assign Upperletter[1431] = 12'b111111111111;
assign Upperletter[1432] = 12'b111111111111;
assign Upperletter[1433] = 12'b000000000000;
assign Upperletter[1434] = 12'b111111111111;
assign Upperletter[1435] = 12'b111111111111;
assign Upperletter[1436] = 12'b111111111111;
assign Upperletter[1437] = 12'b000000000000;
assign Upperletter[1438] = 12'b111111111111;
assign Upperletter[1439] = 12'b111111111111;
assign Upperletter[1440] = 12'b111111111111;
assign Upperletter[1441] = 12'b000000000000;
assign Upperletter[1442] = 12'b111111111111;
assign Upperletter[1443] = 12'b000000000000;
assign Upperletter[1444] = 12'b111111111111;
assign Upperletter[1445] = 12'b000000000000;
assign Upperletter[1446] = 12'b111111111111;
assign Upperletter[1447] = 12'b111111111111;
assign Upperletter[1448] = 12'b111111111111;
assign Upperletter[1449] = 12'b000000000000;
assign Upperletter[1450] = 12'b000000000000;
assign Upperletter[1451] = 12'b111111111111;
assign Upperletter[1452] = 12'b000000000000;
assign Upperletter[1453] = 12'b000000000000;
assign Upperletter[1454] = 12'b111111111111;
assign Upperletter[1455] = 12'b111111111111;
assign Upperletter[1456] = 12'b111111111111;
assign Upperletter[1457] = 12'b000000000000;
assign Upperletter[1458] = 12'b111111111111;
assign Upperletter[1459] = 12'b111111111111;
assign Upperletter[1460] = 12'b111111111111;
assign Upperletter[1461] = 12'b000000000000;
assign Upperletter[1462] = 12'b111111111111;
assign Upperletter[1463] = 12'b111111111111;
assign Upperletter[1464] = 12'b111111111111;
assign Upperletter[1465] = 12'b111111111111;
assign Upperletter[1466] = 12'b111111111111;
assign Upperletter[1467] = 12'b111111111111;
assign Upperletter[1468] = 12'b111111111111;
assign Upperletter[1469] = 12'b111111111111;
assign Upperletter[1470] = 12'b111111111111;
assign Upperletter[1471] = 12'b111111111111;
assign Upperletter[1472] = 12'b111111111111;
assign Upperletter[1473] = 12'b000000000000;
assign Upperletter[1474] = 12'b111111111111;
assign Upperletter[1475] = 12'b111111111111;
assign Upperletter[1476] = 12'b111111111111;
assign Upperletter[1477] = 12'b000000000000;
assign Upperletter[1478] = 12'b111111111111;
assign Upperletter[1479] = 12'b111111111111;
assign Upperletter[1480] = 12'b111111111111;
assign Upperletter[1481] = 12'b000000000000;
assign Upperletter[1482] = 12'b111111111111;
assign Upperletter[1483] = 12'b111111111111;
assign Upperletter[1484] = 12'b111111111111;
assign Upperletter[1485] = 12'b000000000000;
assign Upperletter[1486] = 12'b111111111111;
assign Upperletter[1487] = 12'b111111111111;
assign Upperletter[1488] = 12'b111111111111;
assign Upperletter[1489] = 12'b111111111111;
assign Upperletter[1490] = 12'b000000000000;
assign Upperletter[1491] = 12'b111111111111;
assign Upperletter[1492] = 12'b000000000000;
assign Upperletter[1493] = 12'b111111111111;
assign Upperletter[1494] = 12'b111111111111;
assign Upperletter[1495] = 12'b111111111111;
assign Upperletter[1496] = 12'b111111111111;
assign Upperletter[1497] = 12'b111111111111;
assign Upperletter[1498] = 12'b111111111111;
assign Upperletter[1499] = 12'b000000000000;
assign Upperletter[1500] = 12'b111111111111;
assign Upperletter[1501] = 12'b111111111111;
assign Upperletter[1502] = 12'b111111111111;
assign Upperletter[1503] = 12'b111111111111;
assign Upperletter[1504] = 12'b111111111111;
assign Upperletter[1505] = 12'b111111111111;
assign Upperletter[1506] = 12'b000000000000;
assign Upperletter[1507] = 12'b111111111111;
assign Upperletter[1508] = 12'b000000000000;
assign Upperletter[1509] = 12'b111111111111;
assign Upperletter[1510] = 12'b111111111111;
assign Upperletter[1511] = 12'b111111111111;
assign Upperletter[1512] = 12'b111111111111;
assign Upperletter[1513] = 12'b000000000000;
assign Upperletter[1514] = 12'b111111111111;
assign Upperletter[1515] = 12'b111111111111;
assign Upperletter[1516] = 12'b111111111111;
assign Upperletter[1517] = 12'b000000000000;
assign Upperletter[1518] = 12'b111111111111;
assign Upperletter[1519] = 12'b111111111111;
assign Upperletter[1520] = 12'b111111111111;
assign Upperletter[1521] = 12'b000000000000;
assign Upperletter[1522] = 12'b111111111111;
assign Upperletter[1523] = 12'b111111111111;
assign Upperletter[1524] = 12'b111111111111;
assign Upperletter[1525] = 12'b000000000000;
assign Upperletter[1526] = 12'b111111111111;
assign Upperletter[1527] = 12'b111111111111;
assign Upperletter[1528] = 12'b111111111111;
assign Upperletter[1529] = 12'b111111111111;
assign Upperletter[1530] = 12'b111111111111;
assign Upperletter[1531] = 12'b111111111111;
assign Upperletter[1532] = 12'b111111111111;
assign Upperletter[1533] = 12'b111111111111;
assign Upperletter[1534] = 12'b111111111111;
assign Upperletter[1535] = 12'b111111111111;
assign Upperletter[1536] = 12'b111111111111;
assign Upperletter[1537] = 12'b000000000000;
assign Upperletter[1538] = 12'b111111111111;
assign Upperletter[1539] = 12'b111111111111;
assign Upperletter[1540] = 12'b111111111111;
assign Upperletter[1541] = 12'b000000000000;
assign Upperletter[1542] = 12'b111111111111;
assign Upperletter[1543] = 12'b111111111111;
assign Upperletter[1544] = 12'b111111111111;
assign Upperletter[1545] = 12'b000000000000;
assign Upperletter[1546] = 12'b111111111111;
assign Upperletter[1547] = 12'b111111111111;
assign Upperletter[1548] = 12'b111111111111;
assign Upperletter[1549] = 12'b000000000000;
assign Upperletter[1550] = 12'b111111111111;
assign Upperletter[1551] = 12'b111111111111;
assign Upperletter[1552] = 12'b111111111111;
assign Upperletter[1553] = 12'b111111111111;
assign Upperletter[1554] = 12'b000000000000;
assign Upperletter[1555] = 12'b111111111111;
assign Upperletter[1556] = 12'b000000000000;
assign Upperletter[1557] = 12'b111111111111;
assign Upperletter[1558] = 12'b111111111111;
assign Upperletter[1559] = 12'b111111111111;
assign Upperletter[1560] = 12'b111111111111;
assign Upperletter[1561] = 12'b111111111111;
assign Upperletter[1562] = 12'b111111111111;
assign Upperletter[1563] = 12'b000000000000;
assign Upperletter[1564] = 12'b111111111111;
assign Upperletter[1565] = 12'b111111111111;
assign Upperletter[1566] = 12'b111111111111;
assign Upperletter[1567] = 12'b111111111111;
assign Upperletter[1568] = 12'b111111111111;
assign Upperletter[1569] = 12'b111111111111;
assign Upperletter[1570] = 12'b111111111111;
assign Upperletter[1571] = 12'b000000000000;
assign Upperletter[1572] = 12'b111111111111;
assign Upperletter[1573] = 12'b111111111111;
assign Upperletter[1574] = 12'b111111111111;
assign Upperletter[1575] = 12'b111111111111;
assign Upperletter[1576] = 12'b111111111111;
assign Upperletter[1577] = 12'b111111111111;
assign Upperletter[1578] = 12'b111111111111;
assign Upperletter[1579] = 12'b000000000000;
assign Upperletter[1580] = 12'b111111111111;
assign Upperletter[1581] = 12'b111111111111;
assign Upperletter[1582] = 12'b111111111111;
assign Upperletter[1583] = 12'b111111111111;
assign Upperletter[1584] = 12'b111111111111;
assign Upperletter[1585] = 12'b111111111111;
assign Upperletter[1586] = 12'b111111111111;
assign Upperletter[1587] = 12'b000000000000;
assign Upperletter[1588] = 12'b111111111111;
assign Upperletter[1589] = 12'b111111111111;
assign Upperletter[1590] = 12'b111111111111;
assign Upperletter[1591] = 12'b111111111111;
assign Upperletter[1592] = 12'b111111111111;
assign Upperletter[1593] = 12'b111111111111;
assign Upperletter[1594] = 12'b111111111111;
assign Upperletter[1595] = 12'b111111111111;
assign Upperletter[1596] = 12'b111111111111;
assign Upperletter[1597] = 12'b111111111111;
assign Upperletter[1598] = 12'b111111111111;
assign Upperletter[1599] = 12'b111111111111;
assign Upperletter[1600] = 12'b111111111111;
assign Upperletter[1601] = 12'b000000000000;
assign Upperletter[1602] = 12'b000000000000;
assign Upperletter[1603] = 12'b000000000000;
assign Upperletter[1604] = 12'b000000000000;
assign Upperletter[1605] = 12'b000000000000;
assign Upperletter[1606] = 12'b111111111111;
assign Upperletter[1607] = 12'b111111111111;
assign Upperletter[1608] = 12'b111111111111;
assign Upperletter[1609] = 12'b111111111111;
assign Upperletter[1610] = 12'b111111111111;
assign Upperletter[1611] = 12'b111111111111;
assign Upperletter[1612] = 12'b111111111111;
assign Upperletter[1613] = 12'b000000000000;
assign Upperletter[1614] = 12'b111111111111;
assign Upperletter[1615] = 12'b111111111111;
assign Upperletter[1616] = 12'b111111111111;
assign Upperletter[1617] = 12'b111111111111;
assign Upperletter[1618] = 12'b111111111111;
assign Upperletter[1619] = 12'b111111111111;
assign Upperletter[1620] = 12'b000000000000;
assign Upperletter[1621] = 12'b111111111111;
assign Upperletter[1622] = 12'b111111111111;
assign Upperletter[1623] = 12'b111111111111;
assign Upperletter[1624] = 12'b111111111111;
assign Upperletter[1625] = 12'b111111111111;
assign Upperletter[1626] = 12'b111111111111;
assign Upperletter[1627] = 12'b000000000000;
assign Upperletter[1628] = 12'b111111111111;
assign Upperletter[1629] = 12'b111111111111;
assign Upperletter[1630] = 12'b111111111111;
assign Upperletter[1631] = 12'b111111111111;
assign Upperletter[1632] = 12'b111111111111;
assign Upperletter[1633] = 12'b111111111111;
assign Upperletter[1634] = 12'b000000000000;
assign Upperletter[1635] = 12'b111111111111;
assign Upperletter[1636] = 12'b111111111111;
assign Upperletter[1637] = 12'b111111111111;
assign Upperletter[1638] = 12'b111111111111;
assign Upperletter[1639] = 12'b111111111111;
assign Upperletter[1640] = 12'b111111111111;
assign Upperletter[1641] = 12'b000000000000;
assign Upperletter[1642] = 12'b111111111111;
assign Upperletter[1643] = 12'b111111111111;
assign Upperletter[1644] = 12'b111111111111;
assign Upperletter[1645] = 12'b111111111111;
assign Upperletter[1646] = 12'b111111111111;
assign Upperletter[1647] = 12'b111111111111;
assign Upperletter[1648] = 12'b111111111111;
assign Upperletter[1649] = 12'b000000000000;
assign Upperletter[1650] = 12'b000000000000;
assign Upperletter[1651] = 12'b000000000000;
assign Upperletter[1652] = 12'b000000000000;
assign Upperletter[1653] = 12'b000000000000;
assign Upperletter[1654] = 12'b111111111111;
assign Upperletter[1655] = 12'b111111111111;
assign Upperletter[1656] = 12'b111111111111;
assign Upperletter[1657] = 12'b111111111111;
assign Upperletter[1658] = 12'b111111111111;
assign Upperletter[1659] = 12'b111111111111;
assign Upperletter[1660] = 12'b111111111111;
assign Upperletter[1661] = 12'b111111111111;
assign Upperletter[1662] = 12'b111111111111;
assign Upperletter[1663] = 12'b111111111111;
assign CPM[0] = 12'b111111111111;
assign CPM[1] = 12'b111111111111;
assign CPM[2] = 12'b111111111111;
assign CPM[3] = 12'b111111111111;
assign CPM[4] = 12'b111111111111;
assign CPM[5] = 12'b111111111111;
assign CPM[6] = 12'b111111111111;
assign CPM[7] = 12'b111111111111;
assign CPM[8] = 12'b111111111111;
assign CPM[9] = 12'b111111111111;
assign CPM[10] = 12'b111111111111;
assign CPM[11] = 12'b111111111111;
assign CPM[12] = 12'b111111111111;
assign CPM[13] = 12'b111111111111;
assign CPM[14] = 12'b111111111111;
assign CPM[15] = 12'b111111111111;
assign CPM[16] = 12'b111111111111;
assign CPM[17] = 12'b111111111111;
assign CPM[18] = 12'b111111111111;
assign CPM[19] = 12'b111111111111;
assign CPM[20] = 12'b111111111111;
assign CPM[21] = 12'b111111111111;
assign CPM[22] = 12'b111111111111;
assign CPM[23] = 12'b111111111111;
assign CPM[24] = 12'b111111111111;
assign CPM[25] = 12'b111111111111;
assign CPM[26] = 12'b111111111111;
assign CPM[27] = 12'b111111111111;
assign CPM[28] = 12'b111111111111;
assign CPM[29] = 12'b111111111111;
assign CPM[30] = 12'b111111111111;
assign CPM[31] = 12'b111111111111;
assign CPM[32] = 12'b111111111111;
assign CPM[33] = 12'b111111111111;
assign CPM[34] = 12'b111111111111;
assign CPM[35] = 12'b111111111111;
assign CPM[36] = 12'b111111111111;
assign CPM[37] = 12'b111111111111;
assign CPM[38] = 12'b111111111111;
assign CPM[39] = 12'b111111111111;
assign CPM[40] = 12'b111111111111;
assign CPM[41] = 12'b111111111111;
assign CPM[42] = 12'b111111111111;
assign CPM[43] = 12'b111111111111;
assign CPM[44] = 12'b111111111111;
assign CPM[45] = 12'b111111111111;
assign CPM[46] = 12'b111111111111;
assign CPM[47] = 12'b111111111111;
assign CPM[48] = 12'b111111111111;
assign CPM[49] = 12'b111111111111;
assign CPM[50] = 12'b111111111111;
assign CPM[51] = 12'b111111111111;
assign CPM[52] = 12'b111111111111;
assign CPM[53] = 12'b111111111111;
assign CPM[54] = 12'b111111111111;
assign CPM[55] = 12'b111111111111;
assign CPM[56] = 12'b111111111111;
assign CPM[57] = 12'b111111111111;
assign CPM[58] = 12'b111111111111;
assign CPM[59] = 12'b111111111111;
assign CPM[60] = 12'b111111111111;
assign CPM[61] = 12'b111111111111;
assign CPM[62] = 12'b111111111111;
assign CPM[63] = 12'b111111111111;
assign CPM[64] = 12'b111111111111;
assign CPM[65] = 12'b111111111111;
assign CPM[66] = 12'b111111111111;
assign CPM[67] = 12'b111111111111;
assign CPM[68] = 12'b111111111111;
assign CPM[69] = 12'b111111111111;
assign CPM[70] = 12'b111111111111;
assign CPM[71] = 12'b111111111111;
assign CPM[72] = 12'b111111111111;
assign CPM[73] = 12'b111111111111;
assign CPM[74] = 12'b111111111111;
assign CPM[75] = 12'b111111111111;
assign CPM[76] = 12'b111111111111;
assign CPM[77] = 12'b111111111111;
assign CPM[78] = 12'b111111111111;
assign CPM[79] = 12'b111111111111;
assign CPM[80] = 12'b111111111111;
assign CPM[81] = 12'b111111111111;
assign CPM[82] = 12'b111111111111;
assign CPM[83] = 12'b111111111111;
assign CPM[84] = 12'b111111111111;
assign CPM[85] = 12'b111111111111;
assign CPM[86] = 12'b111111111111;
assign CPM[87] = 12'b111111111111;
assign CPM[88] = 12'b111111111111;
assign CPM[89] = 12'b111111111111;
assign CPM[90] = 12'b111111111111;
assign CPM[91] = 12'b111111111111;
assign CPM[92] = 12'b111111111111;
assign CPM[93] = 12'b111111111111;
assign CPM[94] = 12'b111111111111;
assign CPM[95] = 12'b111111111111;
assign CPM[96] = 12'b111111111111;
assign CPM[97] = 12'b111111111111;
assign CPM[98] = 12'b111111111111;
assign CPM[99] = 12'b111111111111;
assign CPM[100] = 12'b111111111111;
assign CPM[101] = 12'b111111111111;
assign CPM[102] = 12'b111111111111;
assign CPM[103] = 12'b111111111111;
assign CPM[104] = 12'b111111111111;
assign CPM[105] = 12'b111111111111;
assign CPM[106] = 12'b111111111111;
assign CPM[107] = 12'b111111111111;
assign CPM[108] = 12'b111111111111;
assign CPM[109] = 12'b111111111111;
assign CPM[110] = 12'b111111111111;
assign CPM[111] = 12'b111111111111;
assign CPM[112] = 12'b111111111111;
assign CPM[113] = 12'b111111111111;
assign CPM[114] = 12'b111111111111;
assign CPM[115] = 12'b111111111111;
assign CPM[116] = 12'b111111111111;
assign CPM[117] = 12'b111111111111;
assign CPM[118] = 12'b111111111111;
assign CPM[119] = 12'b111111111111;
assign CPM[120] = 12'b111111111111;
assign CPM[121] = 12'b111111111111;
assign CPM[122] = 12'b111111111111;
assign CPM[123] = 12'b111111111111;
assign CPM[124] = 12'b111111111111;
assign CPM[125] = 12'b111111111111;
assign CPM[126] = 12'b111111111111;
assign CPM[127] = 12'b111111111111;
assign CPM[128] = 12'b111111111111;
assign CPM[129] = 12'b111111111111;
assign CPM[130] = 12'b111111111111;
assign CPM[131] = 12'b111111111111;
assign CPM[132] = 12'b111111111111;
assign CPM[133] = 12'b111111111111;
assign CPM[134] = 12'b111111111111;
assign CPM[135] = 12'b111111111111;
assign CPM[136] = 12'b000000000000;
assign CPM[137] = 12'b000000000000;
assign CPM[138] = 12'b000000000000;
assign CPM[139] = 12'b000000000000;
assign CPM[140] = 12'b000000000000;
assign CPM[141] = 12'b000000000000;
assign CPM[142] = 12'b000000000000;
assign CPM[143] = 12'b000000000000;
assign CPM[144] = 12'b000000000000;
assign CPM[145] = 12'b000000000000;
assign CPM[146] = 12'b000000000000;
assign CPM[147] = 12'b000000000000;
assign CPM[148] = 12'b000000000000;
assign CPM[149] = 12'b111111111111;
assign CPM[150] = 12'b111111111111;
assign CPM[151] = 12'b111111111111;
assign CPM[152] = 12'b111111111111;
assign CPM[153] = 12'b111111111111;
assign CPM[154] = 12'b111111111111;
assign CPM[155] = 12'b111111111111;
assign CPM[156] = 12'b111111111111;
assign CPM[157] = 12'b111111111111;
assign CPM[158] = 12'b111111111111;
assign CPM[159] = 12'b111111111111;
assign CPM[160] = 12'b111111111111;
assign CPM[161] = 12'b111111111111;
assign CPM[162] = 12'b111111111111;
assign CPM[163] = 12'b111111111111;
assign CPM[164] = 12'b111111111111;
assign CPM[165] = 12'b111111111111;
assign CPM[166] = 12'b111111111111;
assign CPM[167] = 12'b111111111111;
assign CPM[168] = 12'b000000000000;
assign CPM[169] = 12'b000000000000;
assign CPM[170] = 12'b000000000000;
assign CPM[171] = 12'b000000000000;
assign CPM[172] = 12'b000000000000;
assign CPM[173] = 12'b000000000000;
assign CPM[174] = 12'b000000000000;
assign CPM[175] = 12'b000000000000;
assign CPM[176] = 12'b000000000000;
assign CPM[177] = 12'b000000000000;
assign CPM[178] = 12'b000000000000;
assign CPM[179] = 12'b000000000000;
assign CPM[180] = 12'b000000000000;
assign CPM[181] = 12'b111111111111;
assign CPM[182] = 12'b111111111111;
assign CPM[183] = 12'b111111111111;
assign CPM[184] = 12'b111111111111;
assign CPM[185] = 12'b111111111111;
assign CPM[186] = 12'b111111111111;
assign CPM[187] = 12'b111111111111;
assign CPM[188] = 12'b111111111111;
assign CPM[189] = 12'b111111111111;
assign CPM[190] = 12'b111111111111;
assign CPM[191] = 12'b111111111111;
assign CPM[192] = 12'b111111111111;
assign CPM[193] = 12'b111111111111;
assign CPM[194] = 12'b111111111111;
assign CPM[195] = 12'b111111111111;
assign CPM[196] = 12'b111111111111;
assign CPM[197] = 12'b111111111111;
assign CPM[198] = 12'b111111111111;
assign CPM[199] = 12'b111111111111;
assign CPM[200] = 12'b000000000000;
assign CPM[201] = 12'b000000000000;
assign CPM[202] = 12'b000000000000;
assign CPM[203] = 12'b000000000000;
assign CPM[204] = 12'b000000000000;
assign CPM[205] = 12'b000000000000;
assign CPM[206] = 12'b000000000000;
assign CPM[207] = 12'b000000000000;
assign CPM[208] = 12'b000000000000;
assign CPM[209] = 12'b000000000000;
assign CPM[210] = 12'b000000000000;
assign CPM[211] = 12'b000000000000;
assign CPM[212] = 12'b000000000000;
assign CPM[213] = 12'b111111111111;
assign CPM[214] = 12'b111111111111;
assign CPM[215] = 12'b111111111111;
assign CPM[216] = 12'b111111111111;
assign CPM[217] = 12'b111111111111;
assign CPM[218] = 12'b111111111111;
assign CPM[219] = 12'b111111111111;
assign CPM[220] = 12'b111111111111;
assign CPM[221] = 12'b111111111111;
assign CPM[222] = 12'b111111111111;
assign CPM[223] = 12'b111111111111;
assign CPM[224] = 12'b111111111111;
assign CPM[225] = 12'b111111111111;
assign CPM[226] = 12'b111111111111;
assign CPM[227] = 12'b111111111111;
assign CPM[228] = 12'b111111111111;
assign CPM[229] = 12'b111111111111;
assign CPM[230] = 12'b111111111111;
assign CPM[231] = 12'b111111111111;
assign CPM[232] = 12'b000000000000;
assign CPM[233] = 12'b000000000000;
assign CPM[234] = 12'b000000000000;
assign CPM[235] = 12'b000000000000;
assign CPM[236] = 12'b000000000000;
assign CPM[237] = 12'b000000000000;
assign CPM[238] = 12'b000000000000;
assign CPM[239] = 12'b000000000000;
assign CPM[240] = 12'b000000000000;
assign CPM[241] = 12'b000000000000;
assign CPM[242] = 12'b000000000000;
assign CPM[243] = 12'b000000000000;
assign CPM[244] = 12'b000000000000;
assign CPM[245] = 12'b111111111111;
assign CPM[246] = 12'b111111111111;
assign CPM[247] = 12'b111111111111;
assign CPM[248] = 12'b111111111111;
assign CPM[249] = 12'b111111111111;
assign CPM[250] = 12'b111111111111;
assign CPM[251] = 12'b111111111111;
assign CPM[252] = 12'b111111111111;
assign CPM[253] = 12'b111111111111;
assign CPM[254] = 12'b111111111111;
assign CPM[255] = 12'b111111111111;
assign CPM[256] = 12'b111111111111;
assign CPM[257] = 12'b111111111111;
assign CPM[258] = 12'b111111111111;
assign CPM[259] = 12'b111111111111;
assign CPM[260] = 12'b000000000000;
assign CPM[261] = 12'b000000000000;
assign CPM[262] = 12'b000000000000;
assign CPM[263] = 12'b000000000000;
assign CPM[264] = 12'b111111111111;
assign CPM[265] = 12'b111111111111;
assign CPM[266] = 12'b111111111111;
assign CPM[267] = 12'b111111111111;
assign CPM[268] = 12'b111111111111;
assign CPM[269] = 12'b111111111111;
assign CPM[270] = 12'b111111111111;
assign CPM[271] = 12'b111111111111;
assign CPM[272] = 12'b111111111111;
assign CPM[273] = 12'b111111111111;
assign CPM[274] = 12'b111111111111;
assign CPM[275] = 12'b111111111111;
assign CPM[276] = 12'b111111111111;
assign CPM[277] = 12'b000000000000;
assign CPM[278] = 12'b000000000000;
assign CPM[279] = 12'b000000000000;
assign CPM[280] = 12'b000000000000;
assign CPM[281] = 12'b111111111111;
assign CPM[282] = 12'b111111111111;
assign CPM[283] = 12'b111111111111;
assign CPM[284] = 12'b111111111111;
assign CPM[285] = 12'b111111111111;
assign CPM[286] = 12'b111111111111;
assign CPM[287] = 12'b111111111111;
assign CPM[288] = 12'b111111111111;
assign CPM[289] = 12'b111111111111;
assign CPM[290] = 12'b111111111111;
assign CPM[291] = 12'b111111111111;
assign CPM[292] = 12'b000000000000;
assign CPM[293] = 12'b000000000000;
assign CPM[294] = 12'b000000000000;
assign CPM[295] = 12'b000000000000;
assign CPM[296] = 12'b111111111111;
assign CPM[297] = 12'b111111111111;
assign CPM[298] = 12'b111111111111;
assign CPM[299] = 12'b111111111111;
assign CPM[300] = 12'b111111111111;
assign CPM[301] = 12'b111111111111;
assign CPM[302] = 12'b111111111111;
assign CPM[303] = 12'b111111111111;
assign CPM[304] = 12'b111111111111;
assign CPM[305] = 12'b111111111111;
assign CPM[306] = 12'b111111111111;
assign CPM[307] = 12'b111111111111;
assign CPM[308] = 12'b111111111111;
assign CPM[309] = 12'b000000000000;
assign CPM[310] = 12'b000000000000;
assign CPM[311] = 12'b000000000000;
assign CPM[312] = 12'b000000000000;
assign CPM[313] = 12'b111111111111;
assign CPM[314] = 12'b111111111111;
assign CPM[315] = 12'b111111111111;
assign CPM[316] = 12'b111111111111;
assign CPM[317] = 12'b111111111111;
assign CPM[318] = 12'b111111111111;
assign CPM[319] = 12'b111111111111;
assign CPM[320] = 12'b111111111111;
assign CPM[321] = 12'b111111111111;
assign CPM[322] = 12'b111111111111;
assign CPM[323] = 12'b111111111111;
assign CPM[324] = 12'b000000000000;
assign CPM[325] = 12'b000000000000;
assign CPM[326] = 12'b000000000000;
assign CPM[327] = 12'b000000000000;
assign CPM[328] = 12'b111111111111;
assign CPM[329] = 12'b111111111111;
assign CPM[330] = 12'b111111111111;
assign CPM[331] = 12'b111111111111;
assign CPM[332] = 12'b111111111111;
assign CPM[333] = 12'b111111111111;
assign CPM[334] = 12'b111111111111;
assign CPM[335] = 12'b111111111111;
assign CPM[336] = 12'b111111111111;
assign CPM[337] = 12'b111111111111;
assign CPM[338] = 12'b111111111111;
assign CPM[339] = 12'b111111111111;
assign CPM[340] = 12'b111111111111;
assign CPM[341] = 12'b000000000000;
assign CPM[342] = 12'b000000000000;
assign CPM[343] = 12'b000000000000;
assign CPM[344] = 12'b000000000000;
assign CPM[345] = 12'b111111111111;
assign CPM[346] = 12'b111111111111;
assign CPM[347] = 12'b111111111111;
assign CPM[348] = 12'b111111111111;
assign CPM[349] = 12'b111111111111;
assign CPM[350] = 12'b111111111111;
assign CPM[351] = 12'b111111111111;
assign CPM[352] = 12'b111111111111;
assign CPM[353] = 12'b111111111111;
assign CPM[354] = 12'b111111111111;
assign CPM[355] = 12'b111111111111;
assign CPM[356] = 12'b000000000000;
assign CPM[357] = 12'b000000000000;
assign CPM[358] = 12'b000000000000;
assign CPM[359] = 12'b000000000000;
assign CPM[360] = 12'b111111111111;
assign CPM[361] = 12'b111111111111;
assign CPM[362] = 12'b111111111111;
assign CPM[363] = 12'b111111111111;
assign CPM[364] = 12'b111111111111;
assign CPM[365] = 12'b111111111111;
assign CPM[366] = 12'b111111111111;
assign CPM[367] = 12'b111111111111;
assign CPM[368] = 12'b111111111111;
assign CPM[369] = 12'b111111111111;
assign CPM[370] = 12'b111111111111;
assign CPM[371] = 12'b111111111111;
assign CPM[372] = 12'b111111111111;
assign CPM[373] = 12'b000000000000;
assign CPM[374] = 12'b000000000000;
assign CPM[375] = 12'b000000000000;
assign CPM[376] = 12'b000000000000;
assign CPM[377] = 12'b111111111111;
assign CPM[378] = 12'b111111111111;
assign CPM[379] = 12'b111111111111;
assign CPM[380] = 12'b111111111111;
assign CPM[381] = 12'b111111111111;
assign CPM[382] = 12'b111111111111;
assign CPM[383] = 12'b111111111111;
assign CPM[384] = 12'b111111111111;
assign CPM[385] = 12'b111111111111;
assign CPM[386] = 12'b111111111111;
assign CPM[387] = 12'b111111111111;
assign CPM[388] = 12'b000000000000;
assign CPM[389] = 12'b000000000000;
assign CPM[390] = 12'b000000000000;
assign CPM[391] = 12'b000000000000;
assign CPM[392] = 12'b111111111111;
assign CPM[393] = 12'b111111111111;
assign CPM[394] = 12'b111111111111;
assign CPM[395] = 12'b111111111111;
assign CPM[396] = 12'b111111111111;
assign CPM[397] = 12'b111111111111;
assign CPM[398] = 12'b111111111111;
assign CPM[399] = 12'b111111111111;
assign CPM[400] = 12'b111111111111;
assign CPM[401] = 12'b111111111111;
assign CPM[402] = 12'b111111111111;
assign CPM[403] = 12'b111111111111;
assign CPM[404] = 12'b111111111111;
assign CPM[405] = 12'b111111111111;
assign CPM[406] = 12'b111111111111;
assign CPM[407] = 12'b111111111111;
assign CPM[408] = 12'b111111111111;
assign CPM[409] = 12'b111111111111;
assign CPM[410] = 12'b111111111111;
assign CPM[411] = 12'b111111111111;
assign CPM[412] = 12'b111111111111;
assign CPM[413] = 12'b111111111111;
assign CPM[414] = 12'b111111111111;
assign CPM[415] = 12'b111111111111;
assign CPM[416] = 12'b111111111111;
assign CPM[417] = 12'b111111111111;
assign CPM[418] = 12'b111111111111;
assign CPM[419] = 12'b111111111111;
assign CPM[420] = 12'b000000000000;
assign CPM[421] = 12'b000000000000;
assign CPM[422] = 12'b000000000000;
assign CPM[423] = 12'b000000000000;
assign CPM[424] = 12'b111111111111;
assign CPM[425] = 12'b111111111111;
assign CPM[426] = 12'b111111111111;
assign CPM[427] = 12'b111111111111;
assign CPM[428] = 12'b111111111111;
assign CPM[429] = 12'b111111111111;
assign CPM[430] = 12'b111111111111;
assign CPM[431] = 12'b111111111111;
assign CPM[432] = 12'b111111111111;
assign CPM[433] = 12'b111111111111;
assign CPM[434] = 12'b111111111111;
assign CPM[435] = 12'b111111111111;
assign CPM[436] = 12'b111111111111;
assign CPM[437] = 12'b111111111111;
assign CPM[438] = 12'b111111111111;
assign CPM[439] = 12'b111111111111;
assign CPM[440] = 12'b111111111111;
assign CPM[441] = 12'b111111111111;
assign CPM[442] = 12'b111111111111;
assign CPM[443] = 12'b111111111111;
assign CPM[444] = 12'b111111111111;
assign CPM[445] = 12'b111111111111;
assign CPM[446] = 12'b111111111111;
assign CPM[447] = 12'b111111111111;
assign CPM[448] = 12'b111111111111;
assign CPM[449] = 12'b111111111111;
assign CPM[450] = 12'b111111111111;
assign CPM[451] = 12'b111111111111;
assign CPM[452] = 12'b000000000000;
assign CPM[453] = 12'b000000000000;
assign CPM[454] = 12'b000000000000;
assign CPM[455] = 12'b000000000000;
assign CPM[456] = 12'b111111111111;
assign CPM[457] = 12'b111111111111;
assign CPM[458] = 12'b111111111111;
assign CPM[459] = 12'b111111111111;
assign CPM[460] = 12'b111111111111;
assign CPM[461] = 12'b111111111111;
assign CPM[462] = 12'b111111111111;
assign CPM[463] = 12'b111111111111;
assign CPM[464] = 12'b111111111111;
assign CPM[465] = 12'b111111111111;
assign CPM[466] = 12'b111111111111;
assign CPM[467] = 12'b111111111111;
assign CPM[468] = 12'b111111111111;
assign CPM[469] = 12'b111111111111;
assign CPM[470] = 12'b111111111111;
assign CPM[471] = 12'b111111111111;
assign CPM[472] = 12'b111111111111;
assign CPM[473] = 12'b111111111111;
assign CPM[474] = 12'b111111111111;
assign CPM[475] = 12'b111111111111;
assign CPM[476] = 12'b111111111111;
assign CPM[477] = 12'b111111111111;
assign CPM[478] = 12'b111111111111;
assign CPM[479] = 12'b111111111111;
assign CPM[480] = 12'b111111111111;
assign CPM[481] = 12'b111111111111;
assign CPM[482] = 12'b111111111111;
assign CPM[483] = 12'b111111111111;
assign CPM[484] = 12'b000000000000;
assign CPM[485] = 12'b000000000000;
assign CPM[486] = 12'b000000000000;
assign CPM[487] = 12'b000000000000;
assign CPM[488] = 12'b111111111111;
assign CPM[489] = 12'b111111111111;
assign CPM[490] = 12'b111111111111;
assign CPM[491] = 12'b111111111111;
assign CPM[492] = 12'b111111111111;
assign CPM[493] = 12'b111111111111;
assign CPM[494] = 12'b111111111111;
assign CPM[495] = 12'b111111111111;
assign CPM[496] = 12'b111111111111;
assign CPM[497] = 12'b111111111111;
assign CPM[498] = 12'b111111111111;
assign CPM[499] = 12'b111111111111;
assign CPM[500] = 12'b111111111111;
assign CPM[501] = 12'b111111111111;
assign CPM[502] = 12'b111111111111;
assign CPM[503] = 12'b111111111111;
assign CPM[504] = 12'b111111111111;
assign CPM[505] = 12'b111111111111;
assign CPM[506] = 12'b111111111111;
assign CPM[507] = 12'b111111111111;
assign CPM[508] = 12'b111111111111;
assign CPM[509] = 12'b111111111111;
assign CPM[510] = 12'b111111111111;
assign CPM[511] = 12'b111111111111;
assign CPM[512] = 12'b111111111111;
assign CPM[513] = 12'b111111111111;
assign CPM[514] = 12'b111111111111;
assign CPM[515] = 12'b111111111111;
assign CPM[516] = 12'b000000000000;
assign CPM[517] = 12'b000000000000;
assign CPM[518] = 12'b000000000000;
assign CPM[519] = 12'b000000000000;
assign CPM[520] = 12'b111111111111;
assign CPM[521] = 12'b111111111111;
assign CPM[522] = 12'b111111111111;
assign CPM[523] = 12'b111111111111;
assign CPM[524] = 12'b111111111111;
assign CPM[525] = 12'b111111111111;
assign CPM[526] = 12'b111111111111;
assign CPM[527] = 12'b111111111111;
assign CPM[528] = 12'b111111111111;
assign CPM[529] = 12'b111111111111;
assign CPM[530] = 12'b111111111111;
assign CPM[531] = 12'b111111111111;
assign CPM[532] = 12'b111111111111;
assign CPM[533] = 12'b111111111111;
assign CPM[534] = 12'b111111111111;
assign CPM[535] = 12'b111111111111;
assign CPM[536] = 12'b111111111111;
assign CPM[537] = 12'b111111111111;
assign CPM[538] = 12'b111111111111;
assign CPM[539] = 12'b111111111111;
assign CPM[540] = 12'b111111111111;
assign CPM[541] = 12'b111111111111;
assign CPM[542] = 12'b111111111111;
assign CPM[543] = 12'b111111111111;
assign CPM[544] = 12'b111111111111;
assign CPM[545] = 12'b111111111111;
assign CPM[546] = 12'b111111111111;
assign CPM[547] = 12'b111111111111;
assign CPM[548] = 12'b000000000000;
assign CPM[549] = 12'b000000000000;
assign CPM[550] = 12'b000000000000;
assign CPM[551] = 12'b000000000000;
assign CPM[552] = 12'b111111111111;
assign CPM[553] = 12'b111111111111;
assign CPM[554] = 12'b111111111111;
assign CPM[555] = 12'b111111111111;
assign CPM[556] = 12'b111111111111;
assign CPM[557] = 12'b111111111111;
assign CPM[558] = 12'b111111111111;
assign CPM[559] = 12'b111111111111;
assign CPM[560] = 12'b111111111111;
assign CPM[561] = 12'b111111111111;
assign CPM[562] = 12'b111111111111;
assign CPM[563] = 12'b111111111111;
assign CPM[564] = 12'b111111111111;
assign CPM[565] = 12'b111111111111;
assign CPM[566] = 12'b111111111111;
assign CPM[567] = 12'b111111111111;
assign CPM[568] = 12'b111111111111;
assign CPM[569] = 12'b111111111111;
assign CPM[570] = 12'b111111111111;
assign CPM[571] = 12'b111111111111;
assign CPM[572] = 12'b111111111111;
assign CPM[573] = 12'b111111111111;
assign CPM[574] = 12'b111111111111;
assign CPM[575] = 12'b111111111111;
assign CPM[576] = 12'b111111111111;
assign CPM[577] = 12'b111111111111;
assign CPM[578] = 12'b111111111111;
assign CPM[579] = 12'b111111111111;
assign CPM[580] = 12'b000000000000;
assign CPM[581] = 12'b000000000000;
assign CPM[582] = 12'b000000000000;
assign CPM[583] = 12'b000000000000;
assign CPM[584] = 12'b111111111111;
assign CPM[585] = 12'b111111111111;
assign CPM[586] = 12'b111111111111;
assign CPM[587] = 12'b111111111111;
assign CPM[588] = 12'b111111111111;
assign CPM[589] = 12'b111111111111;
assign CPM[590] = 12'b111111111111;
assign CPM[591] = 12'b111111111111;
assign CPM[592] = 12'b111111111111;
assign CPM[593] = 12'b111111111111;
assign CPM[594] = 12'b111111111111;
assign CPM[595] = 12'b111111111111;
assign CPM[596] = 12'b111111111111;
assign CPM[597] = 12'b111111111111;
assign CPM[598] = 12'b111111111111;
assign CPM[599] = 12'b111111111111;
assign CPM[600] = 12'b111111111111;
assign CPM[601] = 12'b111111111111;
assign CPM[602] = 12'b111111111111;
assign CPM[603] = 12'b111111111111;
assign CPM[604] = 12'b111111111111;
assign CPM[605] = 12'b111111111111;
assign CPM[606] = 12'b111111111111;
assign CPM[607] = 12'b111111111111;
assign CPM[608] = 12'b111111111111;
assign CPM[609] = 12'b111111111111;
assign CPM[610] = 12'b111111111111;
assign CPM[611] = 12'b111111111111;
assign CPM[612] = 12'b000000000000;
assign CPM[613] = 12'b000000000000;
assign CPM[614] = 12'b000000000000;
assign CPM[615] = 12'b000000000000;
assign CPM[616] = 12'b111111111111;
assign CPM[617] = 12'b111111111111;
assign CPM[618] = 12'b111111111111;
assign CPM[619] = 12'b111111111111;
assign CPM[620] = 12'b111111111111;
assign CPM[621] = 12'b111111111111;
assign CPM[622] = 12'b111111111111;
assign CPM[623] = 12'b111111111111;
assign CPM[624] = 12'b111111111111;
assign CPM[625] = 12'b111111111111;
assign CPM[626] = 12'b111111111111;
assign CPM[627] = 12'b111111111111;
assign CPM[628] = 12'b111111111111;
assign CPM[629] = 12'b111111111111;
assign CPM[630] = 12'b111111111111;
assign CPM[631] = 12'b111111111111;
assign CPM[632] = 12'b111111111111;
assign CPM[633] = 12'b111111111111;
assign CPM[634] = 12'b111111111111;
assign CPM[635] = 12'b111111111111;
assign CPM[636] = 12'b111111111111;
assign CPM[637] = 12'b111111111111;
assign CPM[638] = 12'b111111111111;
assign CPM[639] = 12'b111111111111;
assign CPM[640] = 12'b111111111111;
assign CPM[641] = 12'b111111111111;
assign CPM[642] = 12'b111111111111;
assign CPM[643] = 12'b111111111111;
assign CPM[644] = 12'b000000000000;
assign CPM[645] = 12'b000000000000;
assign CPM[646] = 12'b000000000000;
assign CPM[647] = 12'b000000000000;
assign CPM[648] = 12'b111111111111;
assign CPM[649] = 12'b111111111111;
assign CPM[650] = 12'b111111111111;
assign CPM[651] = 12'b111111111111;
assign CPM[652] = 12'b111111111111;
assign CPM[653] = 12'b111111111111;
assign CPM[654] = 12'b111111111111;
assign CPM[655] = 12'b111111111111;
assign CPM[656] = 12'b111111111111;
assign CPM[657] = 12'b111111111111;
assign CPM[658] = 12'b111111111111;
assign CPM[659] = 12'b111111111111;
assign CPM[660] = 12'b111111111111;
assign CPM[661] = 12'b111111111111;
assign CPM[662] = 12'b111111111111;
assign CPM[663] = 12'b111111111111;
assign CPM[664] = 12'b111111111111;
assign CPM[665] = 12'b111111111111;
assign CPM[666] = 12'b111111111111;
assign CPM[667] = 12'b111111111111;
assign CPM[668] = 12'b111111111111;
assign CPM[669] = 12'b111111111111;
assign CPM[670] = 12'b111111111111;
assign CPM[671] = 12'b111111111111;
assign CPM[672] = 12'b111111111111;
assign CPM[673] = 12'b111111111111;
assign CPM[674] = 12'b111111111111;
assign CPM[675] = 12'b111111111111;
assign CPM[676] = 12'b000000000000;
assign CPM[677] = 12'b000000000000;
assign CPM[678] = 12'b000000000000;
assign CPM[679] = 12'b000000000000;
assign CPM[680] = 12'b111111111111;
assign CPM[681] = 12'b111111111111;
assign CPM[682] = 12'b111111111111;
assign CPM[683] = 12'b111111111111;
assign CPM[684] = 12'b111111111111;
assign CPM[685] = 12'b111111111111;
assign CPM[686] = 12'b111111111111;
assign CPM[687] = 12'b111111111111;
assign CPM[688] = 12'b111111111111;
assign CPM[689] = 12'b111111111111;
assign CPM[690] = 12'b111111111111;
assign CPM[691] = 12'b111111111111;
assign CPM[692] = 12'b111111111111;
assign CPM[693] = 12'b000000000000;
assign CPM[694] = 12'b000000000000;
assign CPM[695] = 12'b000000000000;
assign CPM[696] = 12'b000000000000;
assign CPM[697] = 12'b111111111111;
assign CPM[698] = 12'b111111111111;
assign CPM[699] = 12'b111111111111;
assign CPM[700] = 12'b111111111111;
assign CPM[701] = 12'b111111111111;
assign CPM[702] = 12'b111111111111;
assign CPM[703] = 12'b111111111111;
assign CPM[704] = 12'b111111111111;
assign CPM[705] = 12'b111111111111;
assign CPM[706] = 12'b111111111111;
assign CPM[707] = 12'b111111111111;
assign CPM[708] = 12'b000000000000;
assign CPM[709] = 12'b000000000000;
assign CPM[710] = 12'b000000000000;
assign CPM[711] = 12'b000000000000;
assign CPM[712] = 12'b111111111111;
assign CPM[713] = 12'b111111111111;
assign CPM[714] = 12'b111111111111;
assign CPM[715] = 12'b111111111111;
assign CPM[716] = 12'b111111111111;
assign CPM[717] = 12'b111111111111;
assign CPM[718] = 12'b111111111111;
assign CPM[719] = 12'b111111111111;
assign CPM[720] = 12'b111111111111;
assign CPM[721] = 12'b111111111111;
assign CPM[722] = 12'b111111111111;
assign CPM[723] = 12'b111111111111;
assign CPM[724] = 12'b111111111111;
assign CPM[725] = 12'b000000000000;
assign CPM[726] = 12'b000000000000;
assign CPM[727] = 12'b000000000000;
assign CPM[728] = 12'b000000000000;
assign CPM[729] = 12'b111111111111;
assign CPM[730] = 12'b111111111111;
assign CPM[731] = 12'b111111111111;
assign CPM[732] = 12'b111111111111;
assign CPM[733] = 12'b111111111111;
assign CPM[734] = 12'b111111111111;
assign CPM[735] = 12'b111111111111;
assign CPM[736] = 12'b111111111111;
assign CPM[737] = 12'b111111111111;
assign CPM[738] = 12'b111111111111;
assign CPM[739] = 12'b111111111111;
assign CPM[740] = 12'b000000000000;
assign CPM[741] = 12'b000000000000;
assign CPM[742] = 12'b000000000000;
assign CPM[743] = 12'b000000000000;
assign CPM[744] = 12'b111111111111;
assign CPM[745] = 12'b111111111111;
assign CPM[746] = 12'b111111111111;
assign CPM[747] = 12'b111111111111;
assign CPM[748] = 12'b111111111111;
assign CPM[749] = 12'b111111111111;
assign CPM[750] = 12'b111111111111;
assign CPM[751] = 12'b111111111111;
assign CPM[752] = 12'b111111111111;
assign CPM[753] = 12'b111111111111;
assign CPM[754] = 12'b111111111111;
assign CPM[755] = 12'b111111111111;
assign CPM[756] = 12'b111111111111;
assign CPM[757] = 12'b000000000000;
assign CPM[758] = 12'b000000000000;
assign CPM[759] = 12'b000000000000;
assign CPM[760] = 12'b000000000000;
assign CPM[761] = 12'b111111111111;
assign CPM[762] = 12'b111111111111;
assign CPM[763] = 12'b111111111111;
assign CPM[764] = 12'b111111111111;
assign CPM[765] = 12'b111111111111;
assign CPM[766] = 12'b111111111111;
assign CPM[767] = 12'b111111111111;
assign CPM[768] = 12'b111111111111;
assign CPM[769] = 12'b111111111111;
assign CPM[770] = 12'b111111111111;
assign CPM[771] = 12'b111111111111;
assign CPM[772] = 12'b000000000000;
assign CPM[773] = 12'b000000000000;
assign CPM[774] = 12'b000000000000;
assign CPM[775] = 12'b000000000000;
assign CPM[776] = 12'b111111111111;
assign CPM[777] = 12'b111111111111;
assign CPM[778] = 12'b111111111111;
assign CPM[779] = 12'b111111111111;
assign CPM[780] = 12'b111111111111;
assign CPM[781] = 12'b111111111111;
assign CPM[782] = 12'b111111111111;
assign CPM[783] = 12'b111111111111;
assign CPM[784] = 12'b111111111111;
assign CPM[785] = 12'b111111111111;
assign CPM[786] = 12'b111111111111;
assign CPM[787] = 12'b111111111111;
assign CPM[788] = 12'b111111111111;
assign CPM[789] = 12'b000000000000;
assign CPM[790] = 12'b000000000000;
assign CPM[791] = 12'b000000000000;
assign CPM[792] = 12'b000000000000;
assign CPM[793] = 12'b111111111111;
assign CPM[794] = 12'b111111111111;
assign CPM[795] = 12'b111111111111;
assign CPM[796] = 12'b111111111111;
assign CPM[797] = 12'b111111111111;
assign CPM[798] = 12'b111111111111;
assign CPM[799] = 12'b111111111111;
assign CPM[800] = 12'b111111111111;
assign CPM[801] = 12'b111111111111;
assign CPM[802] = 12'b111111111111;
assign CPM[803] = 12'b111111111111;
assign CPM[804] = 12'b111111111111;
assign CPM[805] = 12'b111111111111;
assign CPM[806] = 12'b111111111111;
assign CPM[807] = 12'b111111111111;
assign CPM[808] = 12'b000000000000;
assign CPM[809] = 12'b000000000000;
assign CPM[810] = 12'b000000000000;
assign CPM[811] = 12'b000000000000;
assign CPM[812] = 12'b000000000000;
assign CPM[813] = 12'b000000000000;
assign CPM[814] = 12'b000000000000;
assign CPM[815] = 12'b000000000000;
assign CPM[816] = 12'b000000000000;
assign CPM[817] = 12'b000000000000;
assign CPM[818] = 12'b000000000000;
assign CPM[819] = 12'b000000000000;
assign CPM[820] = 12'b000000000000;
assign CPM[821] = 12'b111111111111;
assign CPM[822] = 12'b111111111111;
assign CPM[823] = 12'b111111111111;
assign CPM[824] = 12'b111111111111;
assign CPM[825] = 12'b111111111111;
assign CPM[826] = 12'b111111111111;
assign CPM[827] = 12'b111111111111;
assign CPM[828] = 12'b111111111111;
assign CPM[829] = 12'b111111111111;
assign CPM[830] = 12'b111111111111;
assign CPM[831] = 12'b111111111111;
assign CPM[832] = 12'b111111111111;
assign CPM[833] = 12'b111111111111;
assign CPM[834] = 12'b111111111111;
assign CPM[835] = 12'b111111111111;
assign CPM[836] = 12'b111111111111;
assign CPM[837] = 12'b111111111111;
assign CPM[838] = 12'b111111111111;
assign CPM[839] = 12'b111111111111;
assign CPM[840] = 12'b000000000000;
assign CPM[841] = 12'b000000000000;
assign CPM[842] = 12'b000000000000;
assign CPM[843] = 12'b000000000000;
assign CPM[844] = 12'b000000000000;
assign CPM[845] = 12'b000000000000;
assign CPM[846] = 12'b000000000000;
assign CPM[847] = 12'b000000000000;
assign CPM[848] = 12'b000000000000;
assign CPM[849] = 12'b000000000000;
assign CPM[850] = 12'b000000000000;
assign CPM[851] = 12'b000000000000;
assign CPM[852] = 12'b000000000000;
assign CPM[853] = 12'b111111111111;
assign CPM[854] = 12'b111111111111;
assign CPM[855] = 12'b111111111111;
assign CPM[856] = 12'b111111111111;
assign CPM[857] = 12'b111111111111;
assign CPM[858] = 12'b111111111111;
assign CPM[859] = 12'b111111111111;
assign CPM[860] = 12'b111111111111;
assign CPM[861] = 12'b111111111111;
assign CPM[862] = 12'b111111111111;
assign CPM[863] = 12'b111111111111;
assign CPM[864] = 12'b111111111111;
assign CPM[865] = 12'b111111111111;
assign CPM[866] = 12'b111111111111;
assign CPM[867] = 12'b111111111111;
assign CPM[868] = 12'b111111111111;
assign CPM[869] = 12'b111111111111;
assign CPM[870] = 12'b111111111111;
assign CPM[871] = 12'b111111111111;
assign CPM[872] = 12'b000000000000;
assign CPM[873] = 12'b000000000000;
assign CPM[874] = 12'b000000000000;
assign CPM[875] = 12'b000000000000;
assign CPM[876] = 12'b000000000000;
assign CPM[877] = 12'b000000000000;
assign CPM[878] = 12'b000000000000;
assign CPM[879] = 12'b000000000000;
assign CPM[880] = 12'b000000000000;
assign CPM[881] = 12'b000000000000;
assign CPM[882] = 12'b000000000000;
assign CPM[883] = 12'b000000000000;
assign CPM[884] = 12'b000000000000;
assign CPM[885] = 12'b111111111111;
assign CPM[886] = 12'b111111111111;
assign CPM[887] = 12'b111111111111;
assign CPM[888] = 12'b111111111111;
assign CPM[889] = 12'b111111111111;
assign CPM[890] = 12'b111111111111;
assign CPM[891] = 12'b111111111111;
assign CPM[892] = 12'b111111111111;
assign CPM[893] = 12'b111111111111;
assign CPM[894] = 12'b111111111111;
assign CPM[895] = 12'b111111111111;
assign CPM[896] = 12'b111111111111;
assign CPM[897] = 12'b111111111111;
assign CPM[898] = 12'b111111111111;
assign CPM[899] = 12'b111111111111;
assign CPM[900] = 12'b111111111111;
assign CPM[901] = 12'b111111111111;
assign CPM[902] = 12'b111111111111;
assign CPM[903] = 12'b111111111111;
assign CPM[904] = 12'b000000000000;
assign CPM[905] = 12'b000000000000;
assign CPM[906] = 12'b000000000000;
assign CPM[907] = 12'b000000000000;
assign CPM[908] = 12'b000000000000;
assign CPM[909] = 12'b000000000000;
assign CPM[910] = 12'b000000000000;
assign CPM[911] = 12'b000000000000;
assign CPM[912] = 12'b000000000000;
assign CPM[913] = 12'b000000000000;
assign CPM[914] = 12'b000000000000;
assign CPM[915] = 12'b000000000000;
assign CPM[916] = 12'b000000000000;
assign CPM[917] = 12'b111111111111;
assign CPM[918] = 12'b111111111111;
assign CPM[919] = 12'b111111111111;
assign CPM[920] = 12'b111111111111;
assign CPM[921] = 12'b111111111111;
assign CPM[922] = 12'b111111111111;
assign CPM[923] = 12'b111111111111;
assign CPM[924] = 12'b111111111111;
assign CPM[925] = 12'b111111111111;
assign CPM[926] = 12'b111111111111;
assign CPM[927] = 12'b111111111111;
assign CPM[928] = 12'b111111111111;
assign CPM[929] = 12'b111111111111;
assign CPM[930] = 12'b111111111111;
assign CPM[931] = 12'b111111111111;
assign CPM[932] = 12'b111111111111;
assign CPM[933] = 12'b111111111111;
assign CPM[934] = 12'b111111111111;
assign CPM[935] = 12'b111111111111;
assign CPM[936] = 12'b111111111111;
assign CPM[937] = 12'b111111111111;
assign CPM[938] = 12'b111111111111;
assign CPM[939] = 12'b111111111111;
assign CPM[940] = 12'b111111111111;
assign CPM[941] = 12'b111111111111;
assign CPM[942] = 12'b111111111111;
assign CPM[943] = 12'b111111111111;
assign CPM[944] = 12'b111111111111;
assign CPM[945] = 12'b111111111111;
assign CPM[946] = 12'b111111111111;
assign CPM[947] = 12'b111111111111;
assign CPM[948] = 12'b111111111111;
assign CPM[949] = 12'b111111111111;
assign CPM[950] = 12'b111111111111;
assign CPM[951] = 12'b111111111111;
assign CPM[952] = 12'b111111111111;
assign CPM[953] = 12'b111111111111;
assign CPM[954] = 12'b111111111111;
assign CPM[955] = 12'b111111111111;
assign CPM[956] = 12'b111111111111;
assign CPM[957] = 12'b111111111111;
assign CPM[958] = 12'b111111111111;
assign CPM[959] = 12'b111111111111;
assign CPM[960] = 12'b111111111111;
assign CPM[961] = 12'b111111111111;
assign CPM[962] = 12'b111111111111;
assign CPM[963] = 12'b111111111111;
assign CPM[964] = 12'b111111111111;
assign CPM[965] = 12'b111111111111;
assign CPM[966] = 12'b111111111111;
assign CPM[967] = 12'b111111111111;
assign CPM[968] = 12'b111111111111;
assign CPM[969] = 12'b111111111111;
assign CPM[970] = 12'b111111111111;
assign CPM[971] = 12'b111111111111;
assign CPM[972] = 12'b111111111111;
assign CPM[973] = 12'b111111111111;
assign CPM[974] = 12'b111111111111;
assign CPM[975] = 12'b111111111111;
assign CPM[976] = 12'b111111111111;
assign CPM[977] = 12'b111111111111;
assign CPM[978] = 12'b111111111111;
assign CPM[979] = 12'b111111111111;
assign CPM[980] = 12'b111111111111;
assign CPM[981] = 12'b111111111111;
assign CPM[982] = 12'b111111111111;
assign CPM[983] = 12'b111111111111;
assign CPM[984] = 12'b111111111111;
assign CPM[985] = 12'b111111111111;
assign CPM[986] = 12'b111111111111;
assign CPM[987] = 12'b111111111111;
assign CPM[988] = 12'b111111111111;
assign CPM[989] = 12'b111111111111;
assign CPM[990] = 12'b111111111111;
assign CPM[991] = 12'b111111111111;
assign CPM[992] = 12'b111111111111;
assign CPM[993] = 12'b111111111111;
assign CPM[994] = 12'b111111111111;
assign CPM[995] = 12'b111111111111;
assign CPM[996] = 12'b111111111111;
assign CPM[997] = 12'b111111111111;
assign CPM[998] = 12'b111111111111;
assign CPM[999] = 12'b111111111111;
assign CPM[1000] = 12'b111111111111;
assign CPM[1001] = 12'b111111111111;
assign CPM[1002] = 12'b111111111111;
assign CPM[1003] = 12'b111111111111;
assign CPM[1004] = 12'b111111111111;
assign CPM[1005] = 12'b111111111111;
assign CPM[1006] = 12'b111111111111;
assign CPM[1007] = 12'b111111111111;
assign CPM[1008] = 12'b111111111111;
assign CPM[1009] = 12'b111111111111;
assign CPM[1010] = 12'b111111111111;
assign CPM[1011] = 12'b111111111111;
assign CPM[1012] = 12'b111111111111;
assign CPM[1013] = 12'b111111111111;
assign CPM[1014] = 12'b111111111111;
assign CPM[1015] = 12'b111111111111;
assign CPM[1016] = 12'b111111111111;
assign CPM[1017] = 12'b111111111111;
assign CPM[1018] = 12'b111111111111;
assign CPM[1019] = 12'b111111111111;
assign CPM[1020] = 12'b111111111111;
assign CPM[1021] = 12'b111111111111;
assign CPM[1022] = 12'b111111111111;
assign CPM[1023] = 12'b111111111111;
assign CPM[1024] = 12'b111111111111;
assign CPM[1025] = 12'b111111111111;
assign CPM[1026] = 12'b111111111111;
assign CPM[1027] = 12'b111111111111;
assign CPM[1028] = 12'b111111111111;
assign CPM[1029] = 12'b111111111111;
assign CPM[1030] = 12'b111111111111;
assign CPM[1031] = 12'b111111111111;
assign CPM[1032] = 12'b111111111111;
assign CPM[1033] = 12'b111111111111;
assign CPM[1034] = 12'b111111111111;
assign CPM[1035] = 12'b111111111111;
assign CPM[1036] = 12'b111111111111;
assign CPM[1037] = 12'b111111111111;
assign CPM[1038] = 12'b111111111111;
assign CPM[1039] = 12'b111111111111;
assign CPM[1040] = 12'b111111111111;
assign CPM[1041] = 12'b111111111111;
assign CPM[1042] = 12'b111111111111;
assign CPM[1043] = 12'b111111111111;
assign CPM[1044] = 12'b111111111111;
assign CPM[1045] = 12'b111111111111;
assign CPM[1046] = 12'b111111111111;
assign CPM[1047] = 12'b111111111111;
assign CPM[1048] = 12'b111111111111;
assign CPM[1049] = 12'b111111111111;
assign CPM[1050] = 12'b111111111111;
assign CPM[1051] = 12'b111111111111;
assign CPM[1052] = 12'b111111111111;
assign CPM[1053] = 12'b111111111111;
assign CPM[1054] = 12'b111111111111;
assign CPM[1055] = 12'b111111111111;
assign CPM[1056] = 12'b111111111111;
assign CPM[1057] = 12'b111111111111;
assign CPM[1058] = 12'b111111111111;
assign CPM[1059] = 12'b111111111111;
assign CPM[1060] = 12'b111111111111;
assign CPM[1061] = 12'b111111111111;
assign CPM[1062] = 12'b111111111111;
assign CPM[1063] = 12'b111111111111;
assign CPM[1064] = 12'b111111111111;
assign CPM[1065] = 12'b111111111111;
assign CPM[1066] = 12'b111111111111;
assign CPM[1067] = 12'b111111111111;
assign CPM[1068] = 12'b111111111111;
assign CPM[1069] = 12'b111111111111;
assign CPM[1070] = 12'b111111111111;
assign CPM[1071] = 12'b111111111111;
assign CPM[1072] = 12'b111111111111;
assign CPM[1073] = 12'b111111111111;
assign CPM[1074] = 12'b111111111111;
assign CPM[1075] = 12'b111111111111;
assign CPM[1076] = 12'b111111111111;
assign CPM[1077] = 12'b111111111111;
assign CPM[1078] = 12'b111111111111;
assign CPM[1079] = 12'b111111111111;
assign CPM[1080] = 12'b111111111111;
assign CPM[1081] = 12'b111111111111;
assign CPM[1082] = 12'b111111111111;
assign CPM[1083] = 12'b111111111111;
assign CPM[1084] = 12'b111111111111;
assign CPM[1085] = 12'b111111111111;
assign CPM[1086] = 12'b111111111111;
assign CPM[1087] = 12'b111111111111;
assign CPM[1088] = 12'b111111111111;
assign CPM[1089] = 12'b111111111111;
assign CPM[1090] = 12'b111111111111;
assign CPM[1091] = 12'b111111111111;
assign CPM[1092] = 12'b111111111111;
assign CPM[1093] = 12'b111111111111;
assign CPM[1094] = 12'b111111111111;
assign CPM[1095] = 12'b111111111111;
assign CPM[1096] = 12'b111111111111;
assign CPM[1097] = 12'b111111111111;
assign CPM[1098] = 12'b111111111111;
assign CPM[1099] = 12'b111111111111;
assign CPM[1100] = 12'b111111111111;
assign CPM[1101] = 12'b111111111111;
assign CPM[1102] = 12'b111111111111;
assign CPM[1103] = 12'b111111111111;
assign CPM[1104] = 12'b111111111111;
assign CPM[1105] = 12'b111111111111;
assign CPM[1106] = 12'b111111111111;
assign CPM[1107] = 12'b111111111111;
assign CPM[1108] = 12'b111111111111;
assign CPM[1109] = 12'b111111111111;
assign CPM[1110] = 12'b111111111111;
assign CPM[1111] = 12'b111111111111;
assign CPM[1112] = 12'b111111111111;
assign CPM[1113] = 12'b111111111111;
assign CPM[1114] = 12'b111111111111;
assign CPM[1115] = 12'b111111111111;
assign CPM[1116] = 12'b111111111111;
assign CPM[1117] = 12'b111111111111;
assign CPM[1118] = 12'b111111111111;
assign CPM[1119] = 12'b111111111111;
assign CPM[1120] = 12'b111111111111;
assign CPM[1121] = 12'b111111111111;
assign CPM[1122] = 12'b111111111111;
assign CPM[1123] = 12'b111111111111;
assign CPM[1124] = 12'b111111111111;
assign CPM[1125] = 12'b000000000000;
assign CPM[1126] = 12'b000000000000;
assign CPM[1127] = 12'b000000000000;
assign CPM[1128] = 12'b000000000000;
assign CPM[1129] = 12'b000000000000;
assign CPM[1130] = 12'b000000000000;
assign CPM[1131] = 12'b000000000000;
assign CPM[1132] = 12'b000000000000;
assign CPM[1133] = 12'b000000000000;
assign CPM[1134] = 12'b000000000000;
assign CPM[1135] = 12'b000000000000;
assign CPM[1136] = 12'b000000000000;
assign CPM[1137] = 12'b000000000000;
assign CPM[1138] = 12'b000000000000;
assign CPM[1139] = 12'b000000000000;
assign CPM[1140] = 12'b000000000000;
assign CPM[1141] = 12'b111111111111;
assign CPM[1142] = 12'b111111111111;
assign CPM[1143] = 12'b111111111111;
assign CPM[1144] = 12'b111111111111;
assign CPM[1145] = 12'b111111111111;
assign CPM[1146] = 12'b111111111111;
assign CPM[1147] = 12'b111111111111;
assign CPM[1148] = 12'b111111111111;
assign CPM[1149] = 12'b111111111111;
assign CPM[1150] = 12'b111111111111;
assign CPM[1151] = 12'b111111111111;
assign CPM[1152] = 12'b111111111111;
assign CPM[1153] = 12'b111111111111;
assign CPM[1154] = 12'b111111111111;
assign CPM[1155] = 12'b111111111111;
assign CPM[1156] = 12'b111111111111;
assign CPM[1157] = 12'b000000000000;
assign CPM[1158] = 12'b000000000000;
assign CPM[1159] = 12'b000000000000;
assign CPM[1160] = 12'b000000000000;
assign CPM[1161] = 12'b000000000000;
assign CPM[1162] = 12'b000000000000;
assign CPM[1163] = 12'b000000000000;
assign CPM[1164] = 12'b000000000000;
assign CPM[1165] = 12'b000000000000;
assign CPM[1166] = 12'b000000000000;
assign CPM[1167] = 12'b000000000000;
assign CPM[1168] = 12'b000000000000;
assign CPM[1169] = 12'b000000000000;
assign CPM[1170] = 12'b000000000000;
assign CPM[1171] = 12'b000000000000;
assign CPM[1172] = 12'b000000000000;
assign CPM[1173] = 12'b111111111111;
assign CPM[1174] = 12'b111111111111;
assign CPM[1175] = 12'b111111111111;
assign CPM[1176] = 12'b111111111111;
assign CPM[1177] = 12'b111111111111;
assign CPM[1178] = 12'b111111111111;
assign CPM[1179] = 12'b111111111111;
assign CPM[1180] = 12'b111111111111;
assign CPM[1181] = 12'b111111111111;
assign CPM[1182] = 12'b111111111111;
assign CPM[1183] = 12'b111111111111;
assign CPM[1184] = 12'b111111111111;
assign CPM[1185] = 12'b111111111111;
assign CPM[1186] = 12'b111111111111;
assign CPM[1187] = 12'b111111111111;
assign CPM[1188] = 12'b111111111111;
assign CPM[1189] = 12'b000000000000;
assign CPM[1190] = 12'b000000000000;
assign CPM[1191] = 12'b000000000000;
assign CPM[1192] = 12'b000000000000;
assign CPM[1193] = 12'b000000000000;
assign CPM[1194] = 12'b000000000000;
assign CPM[1195] = 12'b000000000000;
assign CPM[1196] = 12'b000000000000;
assign CPM[1197] = 12'b000000000000;
assign CPM[1198] = 12'b000000000000;
assign CPM[1199] = 12'b000000000000;
assign CPM[1200] = 12'b000000000000;
assign CPM[1201] = 12'b000000000000;
assign CPM[1202] = 12'b000000000000;
assign CPM[1203] = 12'b000000000000;
assign CPM[1204] = 12'b000000000000;
assign CPM[1205] = 12'b111111111111;
assign CPM[1206] = 12'b111111111111;
assign CPM[1207] = 12'b111111111111;
assign CPM[1208] = 12'b111111111111;
assign CPM[1209] = 12'b111111111111;
assign CPM[1210] = 12'b111111111111;
assign CPM[1211] = 12'b111111111111;
assign CPM[1212] = 12'b111111111111;
assign CPM[1213] = 12'b111111111111;
assign CPM[1214] = 12'b111111111111;
assign CPM[1215] = 12'b111111111111;
assign CPM[1216] = 12'b111111111111;
assign CPM[1217] = 12'b111111111111;
assign CPM[1218] = 12'b111111111111;
assign CPM[1219] = 12'b111111111111;
assign CPM[1220] = 12'b111111111111;
assign CPM[1221] = 12'b000000000000;
assign CPM[1222] = 12'b000000000000;
assign CPM[1223] = 12'b000000000000;
assign CPM[1224] = 12'b000000000000;
assign CPM[1225] = 12'b000000000000;
assign CPM[1226] = 12'b000000000000;
assign CPM[1227] = 12'b000000000000;
assign CPM[1228] = 12'b000000000000;
assign CPM[1229] = 12'b000000000000;
assign CPM[1230] = 12'b000000000000;
assign CPM[1231] = 12'b000000000000;
assign CPM[1232] = 12'b000000000000;
assign CPM[1233] = 12'b000000000000;
assign CPM[1234] = 12'b000000000000;
assign CPM[1235] = 12'b000000000000;
assign CPM[1236] = 12'b000000000000;
assign CPM[1237] = 12'b111111111111;
assign CPM[1238] = 12'b111111111111;
assign CPM[1239] = 12'b111111111111;
assign CPM[1240] = 12'b111111111111;
assign CPM[1241] = 12'b111111111111;
assign CPM[1242] = 12'b111111111111;
assign CPM[1243] = 12'b111111111111;
assign CPM[1244] = 12'b111111111111;
assign CPM[1245] = 12'b111111111111;
assign CPM[1246] = 12'b111111111111;
assign CPM[1247] = 12'b111111111111;
assign CPM[1248] = 12'b111111111111;
assign CPM[1249] = 12'b111111111111;
assign CPM[1250] = 12'b111111111111;
assign CPM[1251] = 12'b111111111111;
assign CPM[1252] = 12'b111111111111;
assign CPM[1253] = 12'b000000000000;
assign CPM[1254] = 12'b000000000000;
assign CPM[1255] = 12'b000000000000;
assign CPM[1256] = 12'b000000000000;
assign CPM[1257] = 12'b111111111111;
assign CPM[1258] = 12'b111111111111;
assign CPM[1259] = 12'b111111111111;
assign CPM[1260] = 12'b111111111111;
assign CPM[1261] = 12'b111111111111;
assign CPM[1262] = 12'b111111111111;
assign CPM[1263] = 12'b111111111111;
assign CPM[1264] = 12'b111111111111;
assign CPM[1265] = 12'b111111111111;
assign CPM[1266] = 12'b111111111111;
assign CPM[1267] = 12'b111111111111;
assign CPM[1268] = 12'b111111111111;
assign CPM[1269] = 12'b000000000000;
assign CPM[1270] = 12'b000000000000;
assign CPM[1271] = 12'b000000000000;
assign CPM[1272] = 12'b000000000000;
assign CPM[1273] = 12'b111111111111;
assign CPM[1274] = 12'b111111111111;
assign CPM[1275] = 12'b111111111111;
assign CPM[1276] = 12'b111111111111;
assign CPM[1277] = 12'b111111111111;
assign CPM[1278] = 12'b111111111111;
assign CPM[1279] = 12'b111111111111;
assign CPM[1280] = 12'b111111111111;
assign CPM[1281] = 12'b111111111111;
assign CPM[1282] = 12'b111111111111;
assign CPM[1283] = 12'b111111111111;
assign CPM[1284] = 12'b111111111111;
assign CPM[1285] = 12'b000000000000;
assign CPM[1286] = 12'b000000000000;
assign CPM[1287] = 12'b000000000000;
assign CPM[1288] = 12'b000000000000;
assign CPM[1289] = 12'b111111111111;
assign CPM[1290] = 12'b111111111111;
assign CPM[1291] = 12'b111111111111;
assign CPM[1292] = 12'b111111111111;
assign CPM[1293] = 12'b111111111111;
assign CPM[1294] = 12'b111111111111;
assign CPM[1295] = 12'b111111111111;
assign CPM[1296] = 12'b111111111111;
assign CPM[1297] = 12'b111111111111;
assign CPM[1298] = 12'b111111111111;
assign CPM[1299] = 12'b111111111111;
assign CPM[1300] = 12'b111111111111;
assign CPM[1301] = 12'b000000000000;
assign CPM[1302] = 12'b000000000000;
assign CPM[1303] = 12'b000000000000;
assign CPM[1304] = 12'b000000000000;
assign CPM[1305] = 12'b111111111111;
assign CPM[1306] = 12'b111111111111;
assign CPM[1307] = 12'b111111111111;
assign CPM[1308] = 12'b111111111111;
assign CPM[1309] = 12'b111111111111;
assign CPM[1310] = 12'b111111111111;
assign CPM[1311] = 12'b111111111111;
assign CPM[1312] = 12'b111111111111;
assign CPM[1313] = 12'b111111111111;
assign CPM[1314] = 12'b111111111111;
assign CPM[1315] = 12'b111111111111;
assign CPM[1316] = 12'b111111111111;
assign CPM[1317] = 12'b000000000000;
assign CPM[1318] = 12'b000000000000;
assign CPM[1319] = 12'b000000000000;
assign CPM[1320] = 12'b000000000000;
assign CPM[1321] = 12'b111111111111;
assign CPM[1322] = 12'b111111111111;
assign CPM[1323] = 12'b111111111111;
assign CPM[1324] = 12'b111111111111;
assign CPM[1325] = 12'b111111111111;
assign CPM[1326] = 12'b111111111111;
assign CPM[1327] = 12'b111111111111;
assign CPM[1328] = 12'b111111111111;
assign CPM[1329] = 12'b111111111111;
assign CPM[1330] = 12'b111111111111;
assign CPM[1331] = 12'b111111111111;
assign CPM[1332] = 12'b111111111111;
assign CPM[1333] = 12'b000000000000;
assign CPM[1334] = 12'b000000000000;
assign CPM[1335] = 12'b000000000000;
assign CPM[1336] = 12'b000000000000;
assign CPM[1337] = 12'b111111111111;
assign CPM[1338] = 12'b111111111111;
assign CPM[1339] = 12'b111111111111;
assign CPM[1340] = 12'b111111111111;
assign CPM[1341] = 12'b111111111111;
assign CPM[1342] = 12'b111111111111;
assign CPM[1343] = 12'b111111111111;
assign CPM[1344] = 12'b111111111111;
assign CPM[1345] = 12'b111111111111;
assign CPM[1346] = 12'b111111111111;
assign CPM[1347] = 12'b111111111111;
assign CPM[1348] = 12'b111111111111;
assign CPM[1349] = 12'b000000000000;
assign CPM[1350] = 12'b000000000000;
assign CPM[1351] = 12'b000000000000;
assign CPM[1352] = 12'b000000000000;
assign CPM[1353] = 12'b111111111111;
assign CPM[1354] = 12'b111111111111;
assign CPM[1355] = 12'b111111111111;
assign CPM[1356] = 12'b111111111111;
assign CPM[1357] = 12'b111111111111;
assign CPM[1358] = 12'b111111111111;
assign CPM[1359] = 12'b111111111111;
assign CPM[1360] = 12'b111111111111;
assign CPM[1361] = 12'b111111111111;
assign CPM[1362] = 12'b111111111111;
assign CPM[1363] = 12'b111111111111;
assign CPM[1364] = 12'b111111111111;
assign CPM[1365] = 12'b000000000000;
assign CPM[1366] = 12'b000000000000;
assign CPM[1367] = 12'b000000000000;
assign CPM[1368] = 12'b000000000000;
assign CPM[1369] = 12'b111111111111;
assign CPM[1370] = 12'b111111111111;
assign CPM[1371] = 12'b111111111111;
assign CPM[1372] = 12'b111111111111;
assign CPM[1373] = 12'b111111111111;
assign CPM[1374] = 12'b111111111111;
assign CPM[1375] = 12'b111111111111;
assign CPM[1376] = 12'b111111111111;
assign CPM[1377] = 12'b111111111111;
assign CPM[1378] = 12'b111111111111;
assign CPM[1379] = 12'b111111111111;
assign CPM[1380] = 12'b111111111111;
assign CPM[1381] = 12'b000000000000;
assign CPM[1382] = 12'b000000000000;
assign CPM[1383] = 12'b000000000000;
assign CPM[1384] = 12'b000000000000;
assign CPM[1385] = 12'b111111111111;
assign CPM[1386] = 12'b111111111111;
assign CPM[1387] = 12'b111111111111;
assign CPM[1388] = 12'b111111111111;
assign CPM[1389] = 12'b111111111111;
assign CPM[1390] = 12'b111111111111;
assign CPM[1391] = 12'b111111111111;
assign CPM[1392] = 12'b111111111111;
assign CPM[1393] = 12'b111111111111;
assign CPM[1394] = 12'b111111111111;
assign CPM[1395] = 12'b111111111111;
assign CPM[1396] = 12'b111111111111;
assign CPM[1397] = 12'b000000000000;
assign CPM[1398] = 12'b000000000000;
assign CPM[1399] = 12'b000000000000;
assign CPM[1400] = 12'b000000000000;
assign CPM[1401] = 12'b111111111111;
assign CPM[1402] = 12'b111111111111;
assign CPM[1403] = 12'b111111111111;
assign CPM[1404] = 12'b111111111111;
assign CPM[1405] = 12'b111111111111;
assign CPM[1406] = 12'b111111111111;
assign CPM[1407] = 12'b111111111111;
assign CPM[1408] = 12'b111111111111;
assign CPM[1409] = 12'b111111111111;
assign CPM[1410] = 12'b111111111111;
assign CPM[1411] = 12'b111111111111;
assign CPM[1412] = 12'b111111111111;
assign CPM[1413] = 12'b000000000000;
assign CPM[1414] = 12'b000000000000;
assign CPM[1415] = 12'b000000000000;
assign CPM[1416] = 12'b000000000000;
assign CPM[1417] = 12'b000000000000;
assign CPM[1418] = 12'b000000000000;
assign CPM[1419] = 12'b000000000000;
assign CPM[1420] = 12'b000000000000;
assign CPM[1421] = 12'b000000000000;
assign CPM[1422] = 12'b000000000000;
assign CPM[1423] = 12'b000000000000;
assign CPM[1424] = 12'b000000000000;
assign CPM[1425] = 12'b000000000000;
assign CPM[1426] = 12'b000000000000;
assign CPM[1427] = 12'b000000000000;
assign CPM[1428] = 12'b000000000000;
assign CPM[1429] = 12'b111111111111;
assign CPM[1430] = 12'b111111111111;
assign CPM[1431] = 12'b111111111111;
assign CPM[1432] = 12'b111111111111;
assign CPM[1433] = 12'b111111111111;
assign CPM[1434] = 12'b111111111111;
assign CPM[1435] = 12'b111111111111;
assign CPM[1436] = 12'b111111111111;
assign CPM[1437] = 12'b111111111111;
assign CPM[1438] = 12'b111111111111;
assign CPM[1439] = 12'b111111111111;
assign CPM[1440] = 12'b111111111111;
assign CPM[1441] = 12'b111111111111;
assign CPM[1442] = 12'b111111111111;
assign CPM[1443] = 12'b111111111111;
assign CPM[1444] = 12'b111111111111;
assign CPM[1445] = 12'b000000000000;
assign CPM[1446] = 12'b000000000000;
assign CPM[1447] = 12'b000000000000;
assign CPM[1448] = 12'b000000000000;
assign CPM[1449] = 12'b000000000000;
assign CPM[1450] = 12'b000000000000;
assign CPM[1451] = 12'b000000000000;
assign CPM[1452] = 12'b000000000000;
assign CPM[1453] = 12'b000000000000;
assign CPM[1454] = 12'b000000000000;
assign CPM[1455] = 12'b000000000000;
assign CPM[1456] = 12'b000000000000;
assign CPM[1457] = 12'b000000000000;
assign CPM[1458] = 12'b000000000000;
assign CPM[1459] = 12'b000000000000;
assign CPM[1460] = 12'b000000000000;
assign CPM[1461] = 12'b111111111111;
assign CPM[1462] = 12'b111111111111;
assign CPM[1463] = 12'b111111111111;
assign CPM[1464] = 12'b111111111111;
assign CPM[1465] = 12'b111111111111;
assign CPM[1466] = 12'b111111111111;
assign CPM[1467] = 12'b111111111111;
assign CPM[1468] = 12'b111111111111;
assign CPM[1469] = 12'b111111111111;
assign CPM[1470] = 12'b111111111111;
assign CPM[1471] = 12'b111111111111;
assign CPM[1472] = 12'b111111111111;
assign CPM[1473] = 12'b111111111111;
assign CPM[1474] = 12'b111111111111;
assign CPM[1475] = 12'b111111111111;
assign CPM[1476] = 12'b111111111111;
assign CPM[1477] = 12'b000000000000;
assign CPM[1478] = 12'b000000000000;
assign CPM[1479] = 12'b000000000000;
assign CPM[1480] = 12'b000000000000;
assign CPM[1481] = 12'b000000000000;
assign CPM[1482] = 12'b000000000000;
assign CPM[1483] = 12'b000000000000;
assign CPM[1484] = 12'b000000000000;
assign CPM[1485] = 12'b000000000000;
assign CPM[1486] = 12'b000000000000;
assign CPM[1487] = 12'b000000000000;
assign CPM[1488] = 12'b000000000000;
assign CPM[1489] = 12'b000000000000;
assign CPM[1490] = 12'b000000000000;
assign CPM[1491] = 12'b000000000000;
assign CPM[1492] = 12'b000000000000;
assign CPM[1493] = 12'b111111111111;
assign CPM[1494] = 12'b111111111111;
assign CPM[1495] = 12'b111111111111;
assign CPM[1496] = 12'b111111111111;
assign CPM[1497] = 12'b111111111111;
assign CPM[1498] = 12'b111111111111;
assign CPM[1499] = 12'b111111111111;
assign CPM[1500] = 12'b111111111111;
assign CPM[1501] = 12'b111111111111;
assign CPM[1502] = 12'b111111111111;
assign CPM[1503] = 12'b111111111111;
assign CPM[1504] = 12'b111111111111;
assign CPM[1505] = 12'b111111111111;
assign CPM[1506] = 12'b111111111111;
assign CPM[1507] = 12'b111111111111;
assign CPM[1508] = 12'b111111111111;
assign CPM[1509] = 12'b000000000000;
assign CPM[1510] = 12'b000000000000;
assign CPM[1511] = 12'b000000000000;
assign CPM[1512] = 12'b000000000000;
assign CPM[1513] = 12'b000000000000;
assign CPM[1514] = 12'b000000000000;
assign CPM[1515] = 12'b000000000000;
assign CPM[1516] = 12'b000000000000;
assign CPM[1517] = 12'b000000000000;
assign CPM[1518] = 12'b000000000000;
assign CPM[1519] = 12'b000000000000;
assign CPM[1520] = 12'b000000000000;
assign CPM[1521] = 12'b000000000000;
assign CPM[1522] = 12'b000000000000;
assign CPM[1523] = 12'b000000000000;
assign CPM[1524] = 12'b000000000000;
assign CPM[1525] = 12'b111111111111;
assign CPM[1526] = 12'b111111111111;
assign CPM[1527] = 12'b111111111111;
assign CPM[1528] = 12'b111111111111;
assign CPM[1529] = 12'b111111111111;
assign CPM[1530] = 12'b111111111111;
assign CPM[1531] = 12'b111111111111;
assign CPM[1532] = 12'b111111111111;
assign CPM[1533] = 12'b111111111111;
assign CPM[1534] = 12'b111111111111;
assign CPM[1535] = 12'b111111111111;
assign CPM[1536] = 12'b111111111111;
assign CPM[1537] = 12'b111111111111;
assign CPM[1538] = 12'b111111111111;
assign CPM[1539] = 12'b111111111111;
assign CPM[1540] = 12'b111111111111;
assign CPM[1541] = 12'b000000000000;
assign CPM[1542] = 12'b000000000000;
assign CPM[1543] = 12'b000000000000;
assign CPM[1544] = 12'b000000000000;
assign CPM[1545] = 12'b111111111111;
assign CPM[1546] = 12'b111111111111;
assign CPM[1547] = 12'b111111111111;
assign CPM[1548] = 12'b111111111111;
assign CPM[1549] = 12'b111111111111;
assign CPM[1550] = 12'b111111111111;
assign CPM[1551] = 12'b111111111111;
assign CPM[1552] = 12'b111111111111;
assign CPM[1553] = 12'b111111111111;
assign CPM[1554] = 12'b111111111111;
assign CPM[1555] = 12'b111111111111;
assign CPM[1556] = 12'b111111111111;
assign CPM[1557] = 12'b111111111111;
assign CPM[1558] = 12'b111111111111;
assign CPM[1559] = 12'b111111111111;
assign CPM[1560] = 12'b111111111111;
assign CPM[1561] = 12'b111111111111;
assign CPM[1562] = 12'b111111111111;
assign CPM[1563] = 12'b111111111111;
assign CPM[1564] = 12'b111111111111;
assign CPM[1565] = 12'b111111111111;
assign CPM[1566] = 12'b111111111111;
assign CPM[1567] = 12'b111111111111;
assign CPM[1568] = 12'b111111111111;
assign CPM[1569] = 12'b111111111111;
assign CPM[1570] = 12'b111111111111;
assign CPM[1571] = 12'b111111111111;
assign CPM[1572] = 12'b111111111111;
assign CPM[1573] = 12'b000000000000;
assign CPM[1574] = 12'b000000000000;
assign CPM[1575] = 12'b000000000000;
assign CPM[1576] = 12'b000000000000;
assign CPM[1577] = 12'b111111111111;
assign CPM[1578] = 12'b111111111111;
assign CPM[1579] = 12'b111111111111;
assign CPM[1580] = 12'b111111111111;
assign CPM[1581] = 12'b111111111111;
assign CPM[1582] = 12'b111111111111;
assign CPM[1583] = 12'b111111111111;
assign CPM[1584] = 12'b111111111111;
assign CPM[1585] = 12'b111111111111;
assign CPM[1586] = 12'b111111111111;
assign CPM[1587] = 12'b111111111111;
assign CPM[1588] = 12'b111111111111;
assign CPM[1589] = 12'b111111111111;
assign CPM[1590] = 12'b111111111111;
assign CPM[1591] = 12'b111111111111;
assign CPM[1592] = 12'b111111111111;
assign CPM[1593] = 12'b111111111111;
assign CPM[1594] = 12'b111111111111;
assign CPM[1595] = 12'b111111111111;
assign CPM[1596] = 12'b111111111111;
assign CPM[1597] = 12'b111111111111;
assign CPM[1598] = 12'b111111111111;
assign CPM[1599] = 12'b111111111111;
assign CPM[1600] = 12'b111111111111;
assign CPM[1601] = 12'b111111111111;
assign CPM[1602] = 12'b111111111111;
assign CPM[1603] = 12'b111111111111;
assign CPM[1604] = 12'b111111111111;
assign CPM[1605] = 12'b000000000000;
assign CPM[1606] = 12'b000000000000;
assign CPM[1607] = 12'b000000000000;
assign CPM[1608] = 12'b000000000000;
assign CPM[1609] = 12'b111111111111;
assign CPM[1610] = 12'b111111111111;
assign CPM[1611] = 12'b111111111111;
assign CPM[1612] = 12'b111111111111;
assign CPM[1613] = 12'b111111111111;
assign CPM[1614] = 12'b111111111111;
assign CPM[1615] = 12'b111111111111;
assign CPM[1616] = 12'b111111111111;
assign CPM[1617] = 12'b111111111111;
assign CPM[1618] = 12'b111111111111;
assign CPM[1619] = 12'b111111111111;
assign CPM[1620] = 12'b111111111111;
assign CPM[1621] = 12'b111111111111;
assign CPM[1622] = 12'b111111111111;
assign CPM[1623] = 12'b111111111111;
assign CPM[1624] = 12'b111111111111;
assign CPM[1625] = 12'b111111111111;
assign CPM[1626] = 12'b111111111111;
assign CPM[1627] = 12'b111111111111;
assign CPM[1628] = 12'b111111111111;
assign CPM[1629] = 12'b111111111111;
assign CPM[1630] = 12'b111111111111;
assign CPM[1631] = 12'b111111111111;
assign CPM[1632] = 12'b111111111111;
assign CPM[1633] = 12'b111111111111;
assign CPM[1634] = 12'b111111111111;
assign CPM[1635] = 12'b111111111111;
assign CPM[1636] = 12'b111111111111;
assign CPM[1637] = 12'b000000000000;
assign CPM[1638] = 12'b000000000000;
assign CPM[1639] = 12'b000000000000;
assign CPM[1640] = 12'b000000000000;
assign CPM[1641] = 12'b111111111111;
assign CPM[1642] = 12'b111111111111;
assign CPM[1643] = 12'b111111111111;
assign CPM[1644] = 12'b111111111111;
assign CPM[1645] = 12'b111111111111;
assign CPM[1646] = 12'b111111111111;
assign CPM[1647] = 12'b111111111111;
assign CPM[1648] = 12'b111111111111;
assign CPM[1649] = 12'b111111111111;
assign CPM[1650] = 12'b111111111111;
assign CPM[1651] = 12'b111111111111;
assign CPM[1652] = 12'b111111111111;
assign CPM[1653] = 12'b111111111111;
assign CPM[1654] = 12'b111111111111;
assign CPM[1655] = 12'b111111111111;
assign CPM[1656] = 12'b111111111111;
assign CPM[1657] = 12'b111111111111;
assign CPM[1658] = 12'b111111111111;
assign CPM[1659] = 12'b111111111111;
assign CPM[1660] = 12'b111111111111;
assign CPM[1661] = 12'b111111111111;
assign CPM[1662] = 12'b111111111111;
assign CPM[1663] = 12'b111111111111;
assign CPM[1664] = 12'b111111111111;
assign CPM[1665] = 12'b111111111111;
assign CPM[1666] = 12'b111111111111;
assign CPM[1667] = 12'b111111111111;
assign CPM[1668] = 12'b111111111111;
assign CPM[1669] = 12'b000000000000;
assign CPM[1670] = 12'b000000000000;
assign CPM[1671] = 12'b000000000000;
assign CPM[1672] = 12'b000000000000;
assign CPM[1673] = 12'b111111111111;
assign CPM[1674] = 12'b111111111111;
assign CPM[1675] = 12'b111111111111;
assign CPM[1676] = 12'b111111111111;
assign CPM[1677] = 12'b111111111111;
assign CPM[1678] = 12'b111111111111;
assign CPM[1679] = 12'b111111111111;
assign CPM[1680] = 12'b111111111111;
assign CPM[1681] = 12'b111111111111;
assign CPM[1682] = 12'b111111111111;
assign CPM[1683] = 12'b111111111111;
assign CPM[1684] = 12'b111111111111;
assign CPM[1685] = 12'b111111111111;
assign CPM[1686] = 12'b111111111111;
assign CPM[1687] = 12'b111111111111;
assign CPM[1688] = 12'b111111111111;
assign CPM[1689] = 12'b111111111111;
assign CPM[1690] = 12'b111111111111;
assign CPM[1691] = 12'b111111111111;
assign CPM[1692] = 12'b111111111111;
assign CPM[1693] = 12'b111111111111;
assign CPM[1694] = 12'b111111111111;
assign CPM[1695] = 12'b111111111111;
assign CPM[1696] = 12'b111111111111;
assign CPM[1697] = 12'b111111111111;
assign CPM[1698] = 12'b111111111111;
assign CPM[1699] = 12'b111111111111;
assign CPM[1700] = 12'b111111111111;
assign CPM[1701] = 12'b000000000000;
assign CPM[1702] = 12'b000000000000;
assign CPM[1703] = 12'b000000000000;
assign CPM[1704] = 12'b000000000000;
assign CPM[1705] = 12'b111111111111;
assign CPM[1706] = 12'b111111111111;
assign CPM[1707] = 12'b111111111111;
assign CPM[1708] = 12'b111111111111;
assign CPM[1709] = 12'b111111111111;
assign CPM[1710] = 12'b111111111111;
assign CPM[1711] = 12'b111111111111;
assign CPM[1712] = 12'b111111111111;
assign CPM[1713] = 12'b111111111111;
assign CPM[1714] = 12'b111111111111;
assign CPM[1715] = 12'b111111111111;
assign CPM[1716] = 12'b111111111111;
assign CPM[1717] = 12'b111111111111;
assign CPM[1718] = 12'b111111111111;
assign CPM[1719] = 12'b111111111111;
assign CPM[1720] = 12'b111111111111;
assign CPM[1721] = 12'b111111111111;
assign CPM[1722] = 12'b111111111111;
assign CPM[1723] = 12'b111111111111;
assign CPM[1724] = 12'b111111111111;
assign CPM[1725] = 12'b111111111111;
assign CPM[1726] = 12'b111111111111;
assign CPM[1727] = 12'b111111111111;
assign CPM[1728] = 12'b111111111111;
assign CPM[1729] = 12'b111111111111;
assign CPM[1730] = 12'b111111111111;
assign CPM[1731] = 12'b111111111111;
assign CPM[1732] = 12'b111111111111;
assign CPM[1733] = 12'b000000000000;
assign CPM[1734] = 12'b000000000000;
assign CPM[1735] = 12'b000000000000;
assign CPM[1736] = 12'b000000000000;
assign CPM[1737] = 12'b111111111111;
assign CPM[1738] = 12'b111111111111;
assign CPM[1739] = 12'b111111111111;
assign CPM[1740] = 12'b111111111111;
assign CPM[1741] = 12'b111111111111;
assign CPM[1742] = 12'b111111111111;
assign CPM[1743] = 12'b111111111111;
assign CPM[1744] = 12'b111111111111;
assign CPM[1745] = 12'b111111111111;
assign CPM[1746] = 12'b111111111111;
assign CPM[1747] = 12'b111111111111;
assign CPM[1748] = 12'b111111111111;
assign CPM[1749] = 12'b111111111111;
assign CPM[1750] = 12'b111111111111;
assign CPM[1751] = 12'b111111111111;
assign CPM[1752] = 12'b111111111111;
assign CPM[1753] = 12'b111111111111;
assign CPM[1754] = 12'b111111111111;
assign CPM[1755] = 12'b111111111111;
assign CPM[1756] = 12'b111111111111;
assign CPM[1757] = 12'b111111111111;
assign CPM[1758] = 12'b111111111111;
assign CPM[1759] = 12'b111111111111;
assign CPM[1760] = 12'b111111111111;
assign CPM[1761] = 12'b111111111111;
assign CPM[1762] = 12'b111111111111;
assign CPM[1763] = 12'b111111111111;
assign CPM[1764] = 12'b111111111111;
assign CPM[1765] = 12'b000000000000;
assign CPM[1766] = 12'b000000000000;
assign CPM[1767] = 12'b000000000000;
assign CPM[1768] = 12'b000000000000;
assign CPM[1769] = 12'b111111111111;
assign CPM[1770] = 12'b111111111111;
assign CPM[1771] = 12'b111111111111;
assign CPM[1772] = 12'b111111111111;
assign CPM[1773] = 12'b111111111111;
assign CPM[1774] = 12'b111111111111;
assign CPM[1775] = 12'b111111111111;
assign CPM[1776] = 12'b111111111111;
assign CPM[1777] = 12'b111111111111;
assign CPM[1778] = 12'b111111111111;
assign CPM[1779] = 12'b111111111111;
assign CPM[1780] = 12'b111111111111;
assign CPM[1781] = 12'b111111111111;
assign CPM[1782] = 12'b111111111111;
assign CPM[1783] = 12'b111111111111;
assign CPM[1784] = 12'b111111111111;
assign CPM[1785] = 12'b111111111111;
assign CPM[1786] = 12'b111111111111;
assign CPM[1787] = 12'b111111111111;
assign CPM[1788] = 12'b111111111111;
assign CPM[1789] = 12'b111111111111;
assign CPM[1790] = 12'b111111111111;
assign CPM[1791] = 12'b111111111111;
assign CPM[1792] = 12'b111111111111;
assign CPM[1793] = 12'b111111111111;
assign CPM[1794] = 12'b111111111111;
assign CPM[1795] = 12'b111111111111;
assign CPM[1796] = 12'b111111111111;
assign CPM[1797] = 12'b000000000000;
assign CPM[1798] = 12'b000000000000;
assign CPM[1799] = 12'b000000000000;
assign CPM[1800] = 12'b000000000000;
assign CPM[1801] = 12'b111111111111;
assign CPM[1802] = 12'b111111111111;
assign CPM[1803] = 12'b111111111111;
assign CPM[1804] = 12'b111111111111;
assign CPM[1805] = 12'b111111111111;
assign CPM[1806] = 12'b111111111111;
assign CPM[1807] = 12'b111111111111;
assign CPM[1808] = 12'b111111111111;
assign CPM[1809] = 12'b111111111111;
assign CPM[1810] = 12'b111111111111;
assign CPM[1811] = 12'b111111111111;
assign CPM[1812] = 12'b111111111111;
assign CPM[1813] = 12'b111111111111;
assign CPM[1814] = 12'b111111111111;
assign CPM[1815] = 12'b111111111111;
assign CPM[1816] = 12'b111111111111;
assign CPM[1817] = 12'b111111111111;
assign CPM[1818] = 12'b111111111111;
assign CPM[1819] = 12'b111111111111;
assign CPM[1820] = 12'b111111111111;
assign CPM[1821] = 12'b111111111111;
assign CPM[1822] = 12'b111111111111;
assign CPM[1823] = 12'b111111111111;
assign CPM[1824] = 12'b111111111111;
assign CPM[1825] = 12'b111111111111;
assign CPM[1826] = 12'b111111111111;
assign CPM[1827] = 12'b111111111111;
assign CPM[1828] = 12'b111111111111;
assign CPM[1829] = 12'b000000000000;
assign CPM[1830] = 12'b000000000000;
assign CPM[1831] = 12'b000000000000;
assign CPM[1832] = 12'b000000000000;
assign CPM[1833] = 12'b111111111111;
assign CPM[1834] = 12'b111111111111;
assign CPM[1835] = 12'b111111111111;
assign CPM[1836] = 12'b111111111111;
assign CPM[1837] = 12'b111111111111;
assign CPM[1838] = 12'b111111111111;
assign CPM[1839] = 12'b111111111111;
assign CPM[1840] = 12'b111111111111;
assign CPM[1841] = 12'b111111111111;
assign CPM[1842] = 12'b111111111111;
assign CPM[1843] = 12'b111111111111;
assign CPM[1844] = 12'b111111111111;
assign CPM[1845] = 12'b111111111111;
assign CPM[1846] = 12'b111111111111;
assign CPM[1847] = 12'b111111111111;
assign CPM[1848] = 12'b111111111111;
assign CPM[1849] = 12'b111111111111;
assign CPM[1850] = 12'b111111111111;
assign CPM[1851] = 12'b111111111111;
assign CPM[1852] = 12'b111111111111;
assign CPM[1853] = 12'b111111111111;
assign CPM[1854] = 12'b111111111111;
assign CPM[1855] = 12'b111111111111;
assign CPM[1856] = 12'b111111111111;
assign CPM[1857] = 12'b111111111111;
assign CPM[1858] = 12'b111111111111;
assign CPM[1859] = 12'b111111111111;
assign CPM[1860] = 12'b111111111111;
assign CPM[1861] = 12'b000000000000;
assign CPM[1862] = 12'b000000000000;
assign CPM[1863] = 12'b000000000000;
assign CPM[1864] = 12'b000000000000;
assign CPM[1865] = 12'b111111111111;
assign CPM[1866] = 12'b111111111111;
assign CPM[1867] = 12'b111111111111;
assign CPM[1868] = 12'b111111111111;
assign CPM[1869] = 12'b111111111111;
assign CPM[1870] = 12'b111111111111;
assign CPM[1871] = 12'b111111111111;
assign CPM[1872] = 12'b111111111111;
assign CPM[1873] = 12'b111111111111;
assign CPM[1874] = 12'b111111111111;
assign CPM[1875] = 12'b111111111111;
assign CPM[1876] = 12'b111111111111;
assign CPM[1877] = 12'b111111111111;
assign CPM[1878] = 12'b111111111111;
assign CPM[1879] = 12'b111111111111;
assign CPM[1880] = 12'b111111111111;
assign CPM[1881] = 12'b111111111111;
assign CPM[1882] = 12'b111111111111;
assign CPM[1883] = 12'b111111111111;
assign CPM[1884] = 12'b111111111111;
assign CPM[1885] = 12'b111111111111;
assign CPM[1886] = 12'b111111111111;
assign CPM[1887] = 12'b111111111111;
assign CPM[1888] = 12'b111111111111;
assign CPM[1889] = 12'b111111111111;
assign CPM[1890] = 12'b111111111111;
assign CPM[1891] = 12'b111111111111;
assign CPM[1892] = 12'b111111111111;
assign CPM[1893] = 12'b000000000000;
assign CPM[1894] = 12'b000000000000;
assign CPM[1895] = 12'b000000000000;
assign CPM[1896] = 12'b000000000000;
assign CPM[1897] = 12'b111111111111;
assign CPM[1898] = 12'b111111111111;
assign CPM[1899] = 12'b111111111111;
assign CPM[1900] = 12'b111111111111;
assign CPM[1901] = 12'b111111111111;
assign CPM[1902] = 12'b111111111111;
assign CPM[1903] = 12'b111111111111;
assign CPM[1904] = 12'b111111111111;
assign CPM[1905] = 12'b111111111111;
assign CPM[1906] = 12'b111111111111;
assign CPM[1907] = 12'b111111111111;
assign CPM[1908] = 12'b111111111111;
assign CPM[1909] = 12'b111111111111;
assign CPM[1910] = 12'b111111111111;
assign CPM[1911] = 12'b111111111111;
assign CPM[1912] = 12'b111111111111;
assign CPM[1913] = 12'b111111111111;
assign CPM[1914] = 12'b111111111111;
assign CPM[1915] = 12'b111111111111;
assign CPM[1916] = 12'b111111111111;
assign CPM[1917] = 12'b111111111111;
assign CPM[1918] = 12'b111111111111;
assign CPM[1919] = 12'b111111111111;
assign CPM[1920] = 12'b111111111111;
assign CPM[1921] = 12'b111111111111;
assign CPM[1922] = 12'b111111111111;
assign CPM[1923] = 12'b111111111111;
assign CPM[1924] = 12'b111111111111;
assign CPM[1925] = 12'b000000000000;
assign CPM[1926] = 12'b000000000000;
assign CPM[1927] = 12'b000000000000;
assign CPM[1928] = 12'b000000000000;
assign CPM[1929] = 12'b111111111111;
assign CPM[1930] = 12'b111111111111;
assign CPM[1931] = 12'b111111111111;
assign CPM[1932] = 12'b111111111111;
assign CPM[1933] = 12'b111111111111;
assign CPM[1934] = 12'b111111111111;
assign CPM[1935] = 12'b111111111111;
assign CPM[1936] = 12'b111111111111;
assign CPM[1937] = 12'b111111111111;
assign CPM[1938] = 12'b111111111111;
assign CPM[1939] = 12'b111111111111;
assign CPM[1940] = 12'b111111111111;
assign CPM[1941] = 12'b111111111111;
assign CPM[1942] = 12'b111111111111;
assign CPM[1943] = 12'b111111111111;
assign CPM[1944] = 12'b111111111111;
assign CPM[1945] = 12'b111111111111;
assign CPM[1946] = 12'b111111111111;
assign CPM[1947] = 12'b111111111111;
assign CPM[1948] = 12'b111111111111;
assign CPM[1949] = 12'b111111111111;
assign CPM[1950] = 12'b111111111111;
assign CPM[1951] = 12'b111111111111;
assign CPM[1952] = 12'b111111111111;
assign CPM[1953] = 12'b111111111111;
assign CPM[1954] = 12'b111111111111;
assign CPM[1955] = 12'b111111111111;
assign CPM[1956] = 12'b111111111111;
assign CPM[1957] = 12'b111111111111;
assign CPM[1958] = 12'b111111111111;
assign CPM[1959] = 12'b111111111111;
assign CPM[1960] = 12'b111111111111;
assign CPM[1961] = 12'b111111111111;
assign CPM[1962] = 12'b111111111111;
assign CPM[1963] = 12'b111111111111;
assign CPM[1964] = 12'b111111111111;
assign CPM[1965] = 12'b111111111111;
assign CPM[1966] = 12'b111111111111;
assign CPM[1967] = 12'b111111111111;
assign CPM[1968] = 12'b111111111111;
assign CPM[1969] = 12'b111111111111;
assign CPM[1970] = 12'b111111111111;
assign CPM[1971] = 12'b111111111111;
assign CPM[1972] = 12'b111111111111;
assign CPM[1973] = 12'b111111111111;
assign CPM[1974] = 12'b111111111111;
assign CPM[1975] = 12'b111111111111;
assign CPM[1976] = 12'b111111111111;
assign CPM[1977] = 12'b111111111111;
assign CPM[1978] = 12'b111111111111;
assign CPM[1979] = 12'b111111111111;
assign CPM[1980] = 12'b111111111111;
assign CPM[1981] = 12'b111111111111;
assign CPM[1982] = 12'b111111111111;
assign CPM[1983] = 12'b111111111111;
assign CPM[1984] = 12'b111111111111;
assign CPM[1985] = 12'b111111111111;
assign CPM[1986] = 12'b111111111111;
assign CPM[1987] = 12'b111111111111;
assign CPM[1988] = 12'b111111111111;
assign CPM[1989] = 12'b111111111111;
assign CPM[1990] = 12'b111111111111;
assign CPM[1991] = 12'b111111111111;
assign CPM[1992] = 12'b111111111111;
assign CPM[1993] = 12'b111111111111;
assign CPM[1994] = 12'b111111111111;
assign CPM[1995] = 12'b111111111111;
assign CPM[1996] = 12'b111111111111;
assign CPM[1997] = 12'b111111111111;
assign CPM[1998] = 12'b111111111111;
assign CPM[1999] = 12'b111111111111;
assign CPM[2000] = 12'b111111111111;
assign CPM[2001] = 12'b111111111111;
assign CPM[2002] = 12'b111111111111;
assign CPM[2003] = 12'b111111111111;
assign CPM[2004] = 12'b111111111111;
assign CPM[2005] = 12'b111111111111;
assign CPM[2006] = 12'b111111111111;
assign CPM[2007] = 12'b111111111111;
assign CPM[2008] = 12'b111111111111;
assign CPM[2009] = 12'b111111111111;
assign CPM[2010] = 12'b111111111111;
assign CPM[2011] = 12'b111111111111;
assign CPM[2012] = 12'b111111111111;
assign CPM[2013] = 12'b111111111111;
assign CPM[2014] = 12'b111111111111;
assign CPM[2015] = 12'b111111111111;
assign CPM[2016] = 12'b111111111111;
assign CPM[2017] = 12'b111111111111;
assign CPM[2018] = 12'b111111111111;
assign CPM[2019] = 12'b111111111111;
assign CPM[2020] = 12'b111111111111;
assign CPM[2021] = 12'b111111111111;
assign CPM[2022] = 12'b111111111111;
assign CPM[2023] = 12'b111111111111;
assign CPM[2024] = 12'b111111111111;
assign CPM[2025] = 12'b111111111111;
assign CPM[2026] = 12'b111111111111;
assign CPM[2027] = 12'b111111111111;
assign CPM[2028] = 12'b111111111111;
assign CPM[2029] = 12'b111111111111;
assign CPM[2030] = 12'b111111111111;
assign CPM[2031] = 12'b111111111111;
assign CPM[2032] = 12'b111111111111;
assign CPM[2033] = 12'b111111111111;
assign CPM[2034] = 12'b111111111111;
assign CPM[2035] = 12'b111111111111;
assign CPM[2036] = 12'b111111111111;
assign CPM[2037] = 12'b111111111111;
assign CPM[2038] = 12'b111111111111;
assign CPM[2039] = 12'b111111111111;
assign CPM[2040] = 12'b111111111111;
assign CPM[2041] = 12'b111111111111;
assign CPM[2042] = 12'b111111111111;
assign CPM[2043] = 12'b111111111111;
assign CPM[2044] = 12'b111111111111;
assign CPM[2045] = 12'b111111111111;
assign CPM[2046] = 12'b111111111111;
assign CPM[2047] = 12'b111111111111;
assign CPM[2048] = 12'b111111111111;
assign CPM[2049] = 12'b111111111111;
assign CPM[2050] = 12'b111111111111;
assign CPM[2051] = 12'b111111111111;
assign CPM[2052] = 12'b111111111111;
assign CPM[2053] = 12'b111111111111;
assign CPM[2054] = 12'b111111111111;
assign CPM[2055] = 12'b111111111111;
assign CPM[2056] = 12'b111111111111;
assign CPM[2057] = 12'b111111111111;
assign CPM[2058] = 12'b111111111111;
assign CPM[2059] = 12'b111111111111;
assign CPM[2060] = 12'b111111111111;
assign CPM[2061] = 12'b111111111111;
assign CPM[2062] = 12'b111111111111;
assign CPM[2063] = 12'b111111111111;
assign CPM[2064] = 12'b111111111111;
assign CPM[2065] = 12'b111111111111;
assign CPM[2066] = 12'b111111111111;
assign CPM[2067] = 12'b111111111111;
assign CPM[2068] = 12'b111111111111;
assign CPM[2069] = 12'b111111111111;
assign CPM[2070] = 12'b111111111111;
assign CPM[2071] = 12'b111111111111;
assign CPM[2072] = 12'b111111111111;
assign CPM[2073] = 12'b111111111111;
assign CPM[2074] = 12'b111111111111;
assign CPM[2075] = 12'b111111111111;
assign CPM[2076] = 12'b111111111111;
assign CPM[2077] = 12'b111111111111;
assign CPM[2078] = 12'b111111111111;
assign CPM[2079] = 12'b111111111111;
assign CPM[2080] = 12'b111111111111;
assign CPM[2081] = 12'b111111111111;
assign CPM[2082] = 12'b111111111111;
assign CPM[2083] = 12'b111111111111;
assign CPM[2084] = 12'b111111111111;
assign CPM[2085] = 12'b111111111111;
assign CPM[2086] = 12'b111111111111;
assign CPM[2087] = 12'b111111111111;
assign CPM[2088] = 12'b111111111111;
assign CPM[2089] = 12'b111111111111;
assign CPM[2090] = 12'b111111111111;
assign CPM[2091] = 12'b111111111111;
assign CPM[2092] = 12'b111111111111;
assign CPM[2093] = 12'b111111111111;
assign CPM[2094] = 12'b111111111111;
assign CPM[2095] = 12'b111111111111;
assign CPM[2096] = 12'b111111111111;
assign CPM[2097] = 12'b111111111111;
assign CPM[2098] = 12'b111111111111;
assign CPM[2099] = 12'b111111111111;
assign CPM[2100] = 12'b111111111111;
assign CPM[2101] = 12'b111111111111;
assign CPM[2102] = 12'b111111111111;
assign CPM[2103] = 12'b111111111111;
assign CPM[2104] = 12'b111111111111;
assign CPM[2105] = 12'b111111111111;
assign CPM[2106] = 12'b111111111111;
assign CPM[2107] = 12'b111111111111;
assign CPM[2108] = 12'b111111111111;
assign CPM[2109] = 12'b111111111111;
assign CPM[2110] = 12'b111111111111;
assign CPM[2111] = 12'b111111111111;
assign CPM[2112] = 12'b111111111111;
assign CPM[2113] = 12'b111111111111;
assign CPM[2114] = 12'b111111111111;
assign CPM[2115] = 12'b111111111111;
assign CPM[2116] = 12'b111111111111;
assign CPM[2117] = 12'b111111111111;
assign CPM[2118] = 12'b111111111111;
assign CPM[2119] = 12'b111111111111;
assign CPM[2120] = 12'b111111111111;
assign CPM[2121] = 12'b111111111111;
assign CPM[2122] = 12'b111111111111;
assign CPM[2123] = 12'b111111111111;
assign CPM[2124] = 12'b111111111111;
assign CPM[2125] = 12'b111111111111;
assign CPM[2126] = 12'b111111111111;
assign CPM[2127] = 12'b111111111111;
assign CPM[2128] = 12'b111111111111;
assign CPM[2129] = 12'b111111111111;
assign CPM[2130] = 12'b111111111111;
assign CPM[2131] = 12'b111111111111;
assign CPM[2132] = 12'b111111111111;
assign CPM[2133] = 12'b111111111111;
assign CPM[2134] = 12'b111111111111;
assign CPM[2135] = 12'b111111111111;
assign CPM[2136] = 12'b111111111111;
assign CPM[2137] = 12'b111111111111;
assign CPM[2138] = 12'b111111111111;
assign CPM[2139] = 12'b111111111111;
assign CPM[2140] = 12'b111111111111;
assign CPM[2141] = 12'b111111111111;
assign CPM[2142] = 12'b111111111111;
assign CPM[2143] = 12'b111111111111;
assign CPM[2144] = 12'b111111111111;
assign CPM[2145] = 12'b111111111111;
assign CPM[2146] = 12'b111111111111;
assign CPM[2147] = 12'b111111111111;
assign CPM[2148] = 12'b000000000000;
assign CPM[2149] = 12'b000000000000;
assign CPM[2150] = 12'b000000000000;
assign CPM[2151] = 12'b000000000000;
assign CPM[2152] = 12'b111111111111;
assign CPM[2153] = 12'b111111111111;
assign CPM[2154] = 12'b111111111111;
assign CPM[2155] = 12'b111111111111;
assign CPM[2156] = 12'b111111111111;
assign CPM[2157] = 12'b111111111111;
assign CPM[2158] = 12'b111111111111;
assign CPM[2159] = 12'b111111111111;
assign CPM[2160] = 12'b111111111111;
assign CPM[2161] = 12'b111111111111;
assign CPM[2162] = 12'b111111111111;
assign CPM[2163] = 12'b111111111111;
assign CPM[2164] = 12'b000000000000;
assign CPM[2165] = 12'b000000000000;
assign CPM[2166] = 12'b000000000000;
assign CPM[2167] = 12'b000000000000;
assign CPM[2168] = 12'b111111111111;
assign CPM[2169] = 12'b111111111111;
assign CPM[2170] = 12'b111111111111;
assign CPM[2171] = 12'b111111111111;
assign CPM[2172] = 12'b111111111111;
assign CPM[2173] = 12'b111111111111;
assign CPM[2174] = 12'b111111111111;
assign CPM[2175] = 12'b111111111111;
assign CPM[2176] = 12'b111111111111;
assign CPM[2177] = 12'b111111111111;
assign CPM[2178] = 12'b111111111111;
assign CPM[2179] = 12'b111111111111;
assign CPM[2180] = 12'b000000000000;
assign CPM[2181] = 12'b000000000000;
assign CPM[2182] = 12'b000000000000;
assign CPM[2183] = 12'b000000000000;
assign CPM[2184] = 12'b111111111111;
assign CPM[2185] = 12'b111111111111;
assign CPM[2186] = 12'b111111111111;
assign CPM[2187] = 12'b111111111111;
assign CPM[2188] = 12'b111111111111;
assign CPM[2189] = 12'b111111111111;
assign CPM[2190] = 12'b111111111111;
assign CPM[2191] = 12'b111111111111;
assign CPM[2192] = 12'b111111111111;
assign CPM[2193] = 12'b111111111111;
assign CPM[2194] = 12'b111111111111;
assign CPM[2195] = 12'b111111111111;
assign CPM[2196] = 12'b000000000000;
assign CPM[2197] = 12'b000000000000;
assign CPM[2198] = 12'b000000000000;
assign CPM[2199] = 12'b000000000000;
assign CPM[2200] = 12'b111111111111;
assign CPM[2201] = 12'b111111111111;
assign CPM[2202] = 12'b111111111111;
assign CPM[2203] = 12'b111111111111;
assign CPM[2204] = 12'b111111111111;
assign CPM[2205] = 12'b111111111111;
assign CPM[2206] = 12'b111111111111;
assign CPM[2207] = 12'b111111111111;
assign CPM[2208] = 12'b111111111111;
assign CPM[2209] = 12'b111111111111;
assign CPM[2210] = 12'b111111111111;
assign CPM[2211] = 12'b111111111111;
assign CPM[2212] = 12'b000000000000;
assign CPM[2213] = 12'b000000000000;
assign CPM[2214] = 12'b000000000000;
assign CPM[2215] = 12'b000000000000;
assign CPM[2216] = 12'b000000000000;
assign CPM[2217] = 12'b000000000000;
assign CPM[2218] = 12'b000000000000;
assign CPM[2219] = 12'b000000000000;
assign CPM[2220] = 12'b111111111111;
assign CPM[2221] = 12'b111111111111;
assign CPM[2222] = 12'b111111111111;
assign CPM[2223] = 12'b111111111111;
assign CPM[2224] = 12'b000000000000;
assign CPM[2225] = 12'b000000000000;
assign CPM[2226] = 12'b000000000000;
assign CPM[2227] = 12'b000000000000;
assign CPM[2228] = 12'b000000000000;
assign CPM[2229] = 12'b000000000000;
assign CPM[2230] = 12'b000000000000;
assign CPM[2231] = 12'b000000000000;
assign CPM[2232] = 12'b111111111111;
assign CPM[2233] = 12'b111111111111;
assign CPM[2234] = 12'b111111111111;
assign CPM[2235] = 12'b111111111111;
assign CPM[2236] = 12'b111111111111;
assign CPM[2237] = 12'b111111111111;
assign CPM[2238] = 12'b111111111111;
assign CPM[2239] = 12'b111111111111;
assign CPM[2240] = 12'b111111111111;
assign CPM[2241] = 12'b111111111111;
assign CPM[2242] = 12'b111111111111;
assign CPM[2243] = 12'b111111111111;
assign CPM[2244] = 12'b000000000000;
assign CPM[2245] = 12'b000000000000;
assign CPM[2246] = 12'b000000000000;
assign CPM[2247] = 12'b000000000000;
assign CPM[2248] = 12'b000000000000;
assign CPM[2249] = 12'b000000000000;
assign CPM[2250] = 12'b000000000000;
assign CPM[2251] = 12'b000000000000;
assign CPM[2252] = 12'b111111111111;
assign CPM[2253] = 12'b111111111111;
assign CPM[2254] = 12'b111111111111;
assign CPM[2255] = 12'b111111111111;
assign CPM[2256] = 12'b000000000000;
assign CPM[2257] = 12'b000000000000;
assign CPM[2258] = 12'b000000000000;
assign CPM[2259] = 12'b000000000000;
assign CPM[2260] = 12'b000000000000;
assign CPM[2261] = 12'b000000000000;
assign CPM[2262] = 12'b000000000000;
assign CPM[2263] = 12'b000000000000;
assign CPM[2264] = 12'b111111111111;
assign CPM[2265] = 12'b111111111111;
assign CPM[2266] = 12'b111111111111;
assign CPM[2267] = 12'b111111111111;
assign CPM[2268] = 12'b111111111111;
assign CPM[2269] = 12'b111111111111;
assign CPM[2270] = 12'b111111111111;
assign CPM[2271] = 12'b111111111111;
assign CPM[2272] = 12'b111111111111;
assign CPM[2273] = 12'b111111111111;
assign CPM[2274] = 12'b111111111111;
assign CPM[2275] = 12'b111111111111;
assign CPM[2276] = 12'b000000000000;
assign CPM[2277] = 12'b000000000000;
assign CPM[2278] = 12'b000000000000;
assign CPM[2279] = 12'b000000000000;
assign CPM[2280] = 12'b000000000000;
assign CPM[2281] = 12'b000000000000;
assign CPM[2282] = 12'b000000000000;
assign CPM[2283] = 12'b000000000000;
assign CPM[2284] = 12'b111111111111;
assign CPM[2285] = 12'b111111111111;
assign CPM[2286] = 12'b111111111111;
assign CPM[2287] = 12'b111111111111;
assign CPM[2288] = 12'b000000000000;
assign CPM[2289] = 12'b000000000000;
assign CPM[2290] = 12'b000000000000;
assign CPM[2291] = 12'b000000000000;
assign CPM[2292] = 12'b000000000000;
assign CPM[2293] = 12'b000000000000;
assign CPM[2294] = 12'b000000000000;
assign CPM[2295] = 12'b000000000000;
assign CPM[2296] = 12'b111111111111;
assign CPM[2297] = 12'b111111111111;
assign CPM[2298] = 12'b111111111111;
assign CPM[2299] = 12'b111111111111;
assign CPM[2300] = 12'b111111111111;
assign CPM[2301] = 12'b111111111111;
assign CPM[2302] = 12'b111111111111;
assign CPM[2303] = 12'b111111111111;
assign CPM[2304] = 12'b111111111111;
assign CPM[2305] = 12'b111111111111;
assign CPM[2306] = 12'b111111111111;
assign CPM[2307] = 12'b111111111111;
assign CPM[2308] = 12'b000000000000;
assign CPM[2309] = 12'b000000000000;
assign CPM[2310] = 12'b000000000000;
assign CPM[2311] = 12'b000000000000;
assign CPM[2312] = 12'b000000000000;
assign CPM[2313] = 12'b000000000000;
assign CPM[2314] = 12'b000000000000;
assign CPM[2315] = 12'b000000000000;
assign CPM[2316] = 12'b111111111111;
assign CPM[2317] = 12'b111111111111;
assign CPM[2318] = 12'b111111111111;
assign CPM[2319] = 12'b111111111111;
assign CPM[2320] = 12'b000000000000;
assign CPM[2321] = 12'b000000000000;
assign CPM[2322] = 12'b000000000000;
assign CPM[2323] = 12'b000000000000;
assign CPM[2324] = 12'b000000000000;
assign CPM[2325] = 12'b000000000000;
assign CPM[2326] = 12'b000000000000;
assign CPM[2327] = 12'b000000000000;
assign CPM[2328] = 12'b111111111111;
assign CPM[2329] = 12'b111111111111;
assign CPM[2330] = 12'b111111111111;
assign CPM[2331] = 12'b111111111111;
assign CPM[2332] = 12'b111111111111;
assign CPM[2333] = 12'b111111111111;
assign CPM[2334] = 12'b111111111111;
assign CPM[2335] = 12'b111111111111;
assign CPM[2336] = 12'b111111111111;
assign CPM[2337] = 12'b111111111111;
assign CPM[2338] = 12'b111111111111;
assign CPM[2339] = 12'b111111111111;
assign CPM[2340] = 12'b000000000000;
assign CPM[2341] = 12'b000000000000;
assign CPM[2342] = 12'b000000000000;
assign CPM[2343] = 12'b000000000000;
assign CPM[2344] = 12'b111111111111;
assign CPM[2345] = 12'b111111111111;
assign CPM[2346] = 12'b111111111111;
assign CPM[2347] = 12'b111111111111;
assign CPM[2348] = 12'b000000000000;
assign CPM[2349] = 12'b000000000000;
assign CPM[2350] = 12'b000000000000;
assign CPM[2351] = 12'b000000000000;
assign CPM[2352] = 12'b111111111111;
assign CPM[2353] = 12'b111111111111;
assign CPM[2354] = 12'b111111111111;
assign CPM[2355] = 12'b111111111111;
assign CPM[2356] = 12'b000000000000;
assign CPM[2357] = 12'b000000000000;
assign CPM[2358] = 12'b000000000000;
assign CPM[2359] = 12'b000000000000;
assign CPM[2360] = 12'b111111111111;
assign CPM[2361] = 12'b111111111111;
assign CPM[2362] = 12'b111111111111;
assign CPM[2363] = 12'b111111111111;
assign CPM[2364] = 12'b111111111111;
assign CPM[2365] = 12'b111111111111;
assign CPM[2366] = 12'b111111111111;
assign CPM[2367] = 12'b111111111111;
assign CPM[2368] = 12'b111111111111;
assign CPM[2369] = 12'b111111111111;
assign CPM[2370] = 12'b111111111111;
assign CPM[2371] = 12'b111111111111;
assign CPM[2372] = 12'b000000000000;
assign CPM[2373] = 12'b000000000000;
assign CPM[2374] = 12'b000000000000;
assign CPM[2375] = 12'b000000000000;
assign CPM[2376] = 12'b111111111111;
assign CPM[2377] = 12'b111111111111;
assign CPM[2378] = 12'b111111111111;
assign CPM[2379] = 12'b111111111111;
assign CPM[2380] = 12'b000000000000;
assign CPM[2381] = 12'b000000000000;
assign CPM[2382] = 12'b000000000000;
assign CPM[2383] = 12'b000000000000;
assign CPM[2384] = 12'b111111111111;
assign CPM[2385] = 12'b111111111111;
assign CPM[2386] = 12'b111111111111;
assign CPM[2387] = 12'b111111111111;
assign CPM[2388] = 12'b000000000000;
assign CPM[2389] = 12'b000000000000;
assign CPM[2390] = 12'b000000000000;
assign CPM[2391] = 12'b000000000000;
assign CPM[2392] = 12'b111111111111;
assign CPM[2393] = 12'b111111111111;
assign CPM[2394] = 12'b111111111111;
assign CPM[2395] = 12'b111111111111;
assign CPM[2396] = 12'b111111111111;
assign CPM[2397] = 12'b111111111111;
assign CPM[2398] = 12'b111111111111;
assign CPM[2399] = 12'b111111111111;
assign CPM[2400] = 12'b111111111111;
assign CPM[2401] = 12'b111111111111;
assign CPM[2402] = 12'b111111111111;
assign CPM[2403] = 12'b111111111111;
assign CPM[2404] = 12'b000000000000;
assign CPM[2405] = 12'b000000000000;
assign CPM[2406] = 12'b000000000000;
assign CPM[2407] = 12'b000000000000;
assign CPM[2408] = 12'b111111111111;
assign CPM[2409] = 12'b111111111111;
assign CPM[2410] = 12'b111111111111;
assign CPM[2411] = 12'b111111111111;
assign CPM[2412] = 12'b000000000000;
assign CPM[2413] = 12'b000000000000;
assign CPM[2414] = 12'b000000000000;
assign CPM[2415] = 12'b000000000000;
assign CPM[2416] = 12'b111111111111;
assign CPM[2417] = 12'b111111111111;
assign CPM[2418] = 12'b111111111111;
assign CPM[2419] = 12'b111111111111;
assign CPM[2420] = 12'b000000000000;
assign CPM[2421] = 12'b000000000000;
assign CPM[2422] = 12'b000000000000;
assign CPM[2423] = 12'b000000000000;
assign CPM[2424] = 12'b111111111111;
assign CPM[2425] = 12'b111111111111;
assign CPM[2426] = 12'b111111111111;
assign CPM[2427] = 12'b111111111111;
assign CPM[2428] = 12'b111111111111;
assign CPM[2429] = 12'b111111111111;
assign CPM[2430] = 12'b111111111111;
assign CPM[2431] = 12'b111111111111;
assign CPM[2432] = 12'b111111111111;
assign CPM[2433] = 12'b111111111111;
assign CPM[2434] = 12'b111111111111;
assign CPM[2435] = 12'b111111111111;
assign CPM[2436] = 12'b000000000000;
assign CPM[2437] = 12'b000000000000;
assign CPM[2438] = 12'b000000000000;
assign CPM[2439] = 12'b000000000000;
assign CPM[2440] = 12'b111111111111;
assign CPM[2441] = 12'b111111111111;
assign CPM[2442] = 12'b111111111111;
assign CPM[2443] = 12'b111111111111;
assign CPM[2444] = 12'b000000000000;
assign CPM[2445] = 12'b000000000000;
assign CPM[2446] = 12'b000000000000;
assign CPM[2447] = 12'b000000000000;
assign CPM[2448] = 12'b111111111111;
assign CPM[2449] = 12'b111111111111;
assign CPM[2450] = 12'b111111111111;
assign CPM[2451] = 12'b111111111111;
assign CPM[2452] = 12'b000000000000;
assign CPM[2453] = 12'b000000000000;
assign CPM[2454] = 12'b000000000000;
assign CPM[2455] = 12'b000000000000;
assign CPM[2456] = 12'b111111111111;
assign CPM[2457] = 12'b111111111111;
assign CPM[2458] = 12'b111111111111;
assign CPM[2459] = 12'b111111111111;
assign CPM[2460] = 12'b111111111111;
assign CPM[2461] = 12'b111111111111;
assign CPM[2462] = 12'b111111111111;
assign CPM[2463] = 12'b111111111111;
assign CPM[2464] = 12'b111111111111;
assign CPM[2465] = 12'b111111111111;
assign CPM[2466] = 12'b111111111111;
assign CPM[2467] = 12'b111111111111;
assign CPM[2468] = 12'b000000000000;
assign CPM[2469] = 12'b000000000000;
assign CPM[2470] = 12'b000000000000;
assign CPM[2471] = 12'b000000000000;
assign CPM[2472] = 12'b111111111111;
assign CPM[2473] = 12'b111111111111;
assign CPM[2474] = 12'b111111111111;
assign CPM[2475] = 12'b111111111111;
assign CPM[2476] = 12'b111111111111;
assign CPM[2477] = 12'b111111111111;
assign CPM[2478] = 12'b111111111111;
assign CPM[2479] = 12'b111111111111;
assign CPM[2480] = 12'b111111111111;
assign CPM[2481] = 12'b111111111111;
assign CPM[2482] = 12'b111111111111;
assign CPM[2483] = 12'b111111111111;
assign CPM[2484] = 12'b000000000000;
assign CPM[2485] = 12'b000000000000;
assign CPM[2486] = 12'b000000000000;
assign CPM[2487] = 12'b000000000000;
assign CPM[2488] = 12'b111111111111;
assign CPM[2489] = 12'b111111111111;
assign CPM[2490] = 12'b111111111111;
assign CPM[2491] = 12'b111111111111;
assign CPM[2492] = 12'b111111111111;
assign CPM[2493] = 12'b111111111111;
assign CPM[2494] = 12'b111111111111;
assign CPM[2495] = 12'b111111111111;
assign CPM[2496] = 12'b111111111111;
assign CPM[2497] = 12'b111111111111;
assign CPM[2498] = 12'b111111111111;
assign CPM[2499] = 12'b111111111111;
assign CPM[2500] = 12'b000000000000;
assign CPM[2501] = 12'b000000000000;
assign CPM[2502] = 12'b000000000000;
assign CPM[2503] = 12'b000000000000;
assign CPM[2504] = 12'b111111111111;
assign CPM[2505] = 12'b111111111111;
assign CPM[2506] = 12'b111111111111;
assign CPM[2507] = 12'b111111111111;
assign CPM[2508] = 12'b111111111111;
assign CPM[2509] = 12'b111111111111;
assign CPM[2510] = 12'b111111111111;
assign CPM[2511] = 12'b111111111111;
assign CPM[2512] = 12'b111111111111;
assign CPM[2513] = 12'b111111111111;
assign CPM[2514] = 12'b111111111111;
assign CPM[2515] = 12'b111111111111;
assign CPM[2516] = 12'b000000000000;
assign CPM[2517] = 12'b000000000000;
assign CPM[2518] = 12'b000000000000;
assign CPM[2519] = 12'b000000000000;
assign CPM[2520] = 12'b111111111111;
assign CPM[2521] = 12'b111111111111;
assign CPM[2522] = 12'b111111111111;
assign CPM[2523] = 12'b111111111111;
assign CPM[2524] = 12'b111111111111;
assign CPM[2525] = 12'b111111111111;
assign CPM[2526] = 12'b111111111111;
assign CPM[2527] = 12'b111111111111;
assign CPM[2528] = 12'b111111111111;
assign CPM[2529] = 12'b111111111111;
assign CPM[2530] = 12'b111111111111;
assign CPM[2531] = 12'b111111111111;
assign CPM[2532] = 12'b000000000000;
assign CPM[2533] = 12'b000000000000;
assign CPM[2534] = 12'b000000000000;
assign CPM[2535] = 12'b000000000000;
assign CPM[2536] = 12'b111111111111;
assign CPM[2537] = 12'b111111111111;
assign CPM[2538] = 12'b111111111111;
assign CPM[2539] = 12'b111111111111;
assign CPM[2540] = 12'b111111111111;
assign CPM[2541] = 12'b111111111111;
assign CPM[2542] = 12'b111111111111;
assign CPM[2543] = 12'b111111111111;
assign CPM[2544] = 12'b111111111111;
assign CPM[2545] = 12'b111111111111;
assign CPM[2546] = 12'b111111111111;
assign CPM[2547] = 12'b111111111111;
assign CPM[2548] = 12'b000000000000;
assign CPM[2549] = 12'b000000000000;
assign CPM[2550] = 12'b000000000000;
assign CPM[2551] = 12'b000000000000;
assign CPM[2552] = 12'b111111111111;
assign CPM[2553] = 12'b111111111111;
assign CPM[2554] = 12'b111111111111;
assign CPM[2555] = 12'b111111111111;
assign CPM[2556] = 12'b111111111111;
assign CPM[2557] = 12'b111111111111;
assign CPM[2558] = 12'b111111111111;
assign CPM[2559] = 12'b111111111111;
assign CPM[2560] = 12'b111111111111;
assign CPM[2561] = 12'b111111111111;
assign CPM[2562] = 12'b111111111111;
assign CPM[2563] = 12'b111111111111;
assign CPM[2564] = 12'b000000000000;
assign CPM[2565] = 12'b000000000000;
assign CPM[2566] = 12'b000000000000;
assign CPM[2567] = 12'b000000000000;
assign CPM[2568] = 12'b111111111111;
assign CPM[2569] = 12'b111111111111;
assign CPM[2570] = 12'b111111111111;
assign CPM[2571] = 12'b111111111111;
assign CPM[2572] = 12'b111111111111;
assign CPM[2573] = 12'b111111111111;
assign CPM[2574] = 12'b111111111111;
assign CPM[2575] = 12'b111111111111;
assign CPM[2576] = 12'b111111111111;
assign CPM[2577] = 12'b111111111111;
assign CPM[2578] = 12'b111111111111;
assign CPM[2579] = 12'b111111111111;
assign CPM[2580] = 12'b000000000000;
assign CPM[2581] = 12'b000000000000;
assign CPM[2582] = 12'b000000000000;
assign CPM[2583] = 12'b000000000000;
assign CPM[2584] = 12'b111111111111;
assign CPM[2585] = 12'b111111111111;
assign CPM[2586] = 12'b111111111111;
assign CPM[2587] = 12'b111111111111;
assign CPM[2588] = 12'b111111111111;
assign CPM[2589] = 12'b111111111111;
assign CPM[2590] = 12'b111111111111;
assign CPM[2591] = 12'b111111111111;
assign CPM[2592] = 12'b111111111111;
assign CPM[2593] = 12'b111111111111;
assign CPM[2594] = 12'b111111111111;
assign CPM[2595] = 12'b111111111111;
assign CPM[2596] = 12'b000000000000;
assign CPM[2597] = 12'b000000000000;
assign CPM[2598] = 12'b000000000000;
assign CPM[2599] = 12'b000000000000;
assign CPM[2600] = 12'b111111111111;
assign CPM[2601] = 12'b111111111111;
assign CPM[2602] = 12'b111111111111;
assign CPM[2603] = 12'b111111111111;
assign CPM[2604] = 12'b111111111111;
assign CPM[2605] = 12'b111111111111;
assign CPM[2606] = 12'b111111111111;
assign CPM[2607] = 12'b111111111111;
assign CPM[2608] = 12'b111111111111;
assign CPM[2609] = 12'b111111111111;
assign CPM[2610] = 12'b111111111111;
assign CPM[2611] = 12'b111111111111;
assign CPM[2612] = 12'b000000000000;
assign CPM[2613] = 12'b000000000000;
assign CPM[2614] = 12'b000000000000;
assign CPM[2615] = 12'b000000000000;
assign CPM[2616] = 12'b111111111111;
assign CPM[2617] = 12'b111111111111;
assign CPM[2618] = 12'b111111111111;
assign CPM[2619] = 12'b111111111111;
assign CPM[2620] = 12'b111111111111;
assign CPM[2621] = 12'b111111111111;
assign CPM[2622] = 12'b111111111111;
assign CPM[2623] = 12'b111111111111;
assign CPM[2624] = 12'b111111111111;
assign CPM[2625] = 12'b111111111111;
assign CPM[2626] = 12'b111111111111;
assign CPM[2627] = 12'b111111111111;
assign CPM[2628] = 12'b000000000000;
assign CPM[2629] = 12'b000000000000;
assign CPM[2630] = 12'b000000000000;
assign CPM[2631] = 12'b000000000000;
assign CPM[2632] = 12'b111111111111;
assign CPM[2633] = 12'b111111111111;
assign CPM[2634] = 12'b111111111111;
assign CPM[2635] = 12'b111111111111;
assign CPM[2636] = 12'b111111111111;
assign CPM[2637] = 12'b111111111111;
assign CPM[2638] = 12'b111111111111;
assign CPM[2639] = 12'b111111111111;
assign CPM[2640] = 12'b111111111111;
assign CPM[2641] = 12'b111111111111;
assign CPM[2642] = 12'b111111111111;
assign CPM[2643] = 12'b111111111111;
assign CPM[2644] = 12'b000000000000;
assign CPM[2645] = 12'b000000000000;
assign CPM[2646] = 12'b000000000000;
assign CPM[2647] = 12'b000000000000;
assign CPM[2648] = 12'b111111111111;
assign CPM[2649] = 12'b111111111111;
assign CPM[2650] = 12'b111111111111;
assign CPM[2651] = 12'b111111111111;
assign CPM[2652] = 12'b111111111111;
assign CPM[2653] = 12'b111111111111;
assign CPM[2654] = 12'b111111111111;
assign CPM[2655] = 12'b111111111111;
assign CPM[2656] = 12'b111111111111;
assign CPM[2657] = 12'b111111111111;
assign CPM[2658] = 12'b111111111111;
assign CPM[2659] = 12'b111111111111;
assign CPM[2660] = 12'b000000000000;
assign CPM[2661] = 12'b000000000000;
assign CPM[2662] = 12'b000000000000;
assign CPM[2663] = 12'b000000000000;
assign CPM[2664] = 12'b111111111111;
assign CPM[2665] = 12'b111111111111;
assign CPM[2666] = 12'b111111111111;
assign CPM[2667] = 12'b111111111111;
assign CPM[2668] = 12'b111111111111;
assign CPM[2669] = 12'b111111111111;
assign CPM[2670] = 12'b111111111111;
assign CPM[2671] = 12'b111111111111;
assign CPM[2672] = 12'b111111111111;
assign CPM[2673] = 12'b111111111111;
assign CPM[2674] = 12'b111111111111;
assign CPM[2675] = 12'b111111111111;
assign CPM[2676] = 12'b000000000000;
assign CPM[2677] = 12'b000000000000;
assign CPM[2678] = 12'b000000000000;
assign CPM[2679] = 12'b000000000000;
assign CPM[2680] = 12'b111111111111;
assign CPM[2681] = 12'b111111111111;
assign CPM[2682] = 12'b111111111111;
assign CPM[2683] = 12'b111111111111;
assign CPM[2684] = 12'b111111111111;
assign CPM[2685] = 12'b111111111111;
assign CPM[2686] = 12'b111111111111;
assign CPM[2687] = 12'b111111111111;
assign CPM[2688] = 12'b111111111111;
assign CPM[2689] = 12'b111111111111;
assign CPM[2690] = 12'b111111111111;
assign CPM[2691] = 12'b111111111111;
assign CPM[2692] = 12'b000000000000;
assign CPM[2693] = 12'b000000000000;
assign CPM[2694] = 12'b000000000000;
assign CPM[2695] = 12'b000000000000;
assign CPM[2696] = 12'b111111111111;
assign CPM[2697] = 12'b111111111111;
assign CPM[2698] = 12'b111111111111;
assign CPM[2699] = 12'b111111111111;
assign CPM[2700] = 12'b111111111111;
assign CPM[2701] = 12'b111111111111;
assign CPM[2702] = 12'b111111111111;
assign CPM[2703] = 12'b111111111111;
assign CPM[2704] = 12'b111111111111;
assign CPM[2705] = 12'b111111111111;
assign CPM[2706] = 12'b111111111111;
assign CPM[2707] = 12'b111111111111;
assign CPM[2708] = 12'b000000000000;
assign CPM[2709] = 12'b000000000000;
assign CPM[2710] = 12'b000000000000;
assign CPM[2711] = 12'b000000000000;
assign CPM[2712] = 12'b111111111111;
assign CPM[2713] = 12'b111111111111;
assign CPM[2714] = 12'b111111111111;
assign CPM[2715] = 12'b111111111111;
assign CPM[2716] = 12'b111111111111;
assign CPM[2717] = 12'b111111111111;
assign CPM[2718] = 12'b111111111111;
assign CPM[2719] = 12'b111111111111;
assign CPM[2720] = 12'b111111111111;
assign CPM[2721] = 12'b111111111111;
assign CPM[2722] = 12'b111111111111;
assign CPM[2723] = 12'b111111111111;
assign CPM[2724] = 12'b000000000000;
assign CPM[2725] = 12'b000000000000;
assign CPM[2726] = 12'b000000000000;
assign CPM[2727] = 12'b000000000000;
assign CPM[2728] = 12'b111111111111;
assign CPM[2729] = 12'b111111111111;
assign CPM[2730] = 12'b111111111111;
assign CPM[2731] = 12'b111111111111;
assign CPM[2732] = 12'b111111111111;
assign CPM[2733] = 12'b111111111111;
assign CPM[2734] = 12'b111111111111;
assign CPM[2735] = 12'b111111111111;
assign CPM[2736] = 12'b111111111111;
assign CPM[2737] = 12'b111111111111;
assign CPM[2738] = 12'b111111111111;
assign CPM[2739] = 12'b111111111111;
assign CPM[2740] = 12'b000000000000;
assign CPM[2741] = 12'b000000000000;
assign CPM[2742] = 12'b000000000000;
assign CPM[2743] = 12'b000000000000;
assign CPM[2744] = 12'b111111111111;
assign CPM[2745] = 12'b111111111111;
assign CPM[2746] = 12'b111111111111;
assign CPM[2747] = 12'b111111111111;
assign CPM[2748] = 12'b111111111111;
assign CPM[2749] = 12'b111111111111;
assign CPM[2750] = 12'b111111111111;
assign CPM[2751] = 12'b111111111111;
assign CPM[2752] = 12'b111111111111;
assign CPM[2753] = 12'b111111111111;
assign CPM[2754] = 12'b111111111111;
assign CPM[2755] = 12'b111111111111;
assign CPM[2756] = 12'b000000000000;
assign CPM[2757] = 12'b000000000000;
assign CPM[2758] = 12'b000000000000;
assign CPM[2759] = 12'b000000000000;
assign CPM[2760] = 12'b111111111111;
assign CPM[2761] = 12'b111111111111;
assign CPM[2762] = 12'b111111111111;
assign CPM[2763] = 12'b111111111111;
assign CPM[2764] = 12'b111111111111;
assign CPM[2765] = 12'b111111111111;
assign CPM[2766] = 12'b111111111111;
assign CPM[2767] = 12'b111111111111;
assign CPM[2768] = 12'b111111111111;
assign CPM[2769] = 12'b111111111111;
assign CPM[2770] = 12'b111111111111;
assign CPM[2771] = 12'b111111111111;
assign CPM[2772] = 12'b000000000000;
assign CPM[2773] = 12'b000000000000;
assign CPM[2774] = 12'b000000000000;
assign CPM[2775] = 12'b000000000000;
assign CPM[2776] = 12'b111111111111;
assign CPM[2777] = 12'b111111111111;
assign CPM[2778] = 12'b111111111111;
assign CPM[2779] = 12'b111111111111;
assign CPM[2780] = 12'b111111111111;
assign CPM[2781] = 12'b111111111111;
assign CPM[2782] = 12'b111111111111;
assign CPM[2783] = 12'b111111111111;
assign CPM[2784] = 12'b111111111111;
assign CPM[2785] = 12'b111111111111;
assign CPM[2786] = 12'b111111111111;
assign CPM[2787] = 12'b111111111111;
assign CPM[2788] = 12'b000000000000;
assign CPM[2789] = 12'b000000000000;
assign CPM[2790] = 12'b000000000000;
assign CPM[2791] = 12'b000000000000;
assign CPM[2792] = 12'b111111111111;
assign CPM[2793] = 12'b111111111111;
assign CPM[2794] = 12'b111111111111;
assign CPM[2795] = 12'b111111111111;
assign CPM[2796] = 12'b111111111111;
assign CPM[2797] = 12'b111111111111;
assign CPM[2798] = 12'b111111111111;
assign CPM[2799] = 12'b111111111111;
assign CPM[2800] = 12'b111111111111;
assign CPM[2801] = 12'b111111111111;
assign CPM[2802] = 12'b111111111111;
assign CPM[2803] = 12'b111111111111;
assign CPM[2804] = 12'b000000000000;
assign CPM[2805] = 12'b000000000000;
assign CPM[2806] = 12'b000000000000;
assign CPM[2807] = 12'b000000000000;
assign CPM[2808] = 12'b111111111111;
assign CPM[2809] = 12'b111111111111;
assign CPM[2810] = 12'b111111111111;
assign CPM[2811] = 12'b111111111111;
assign CPM[2812] = 12'b111111111111;
assign CPM[2813] = 12'b111111111111;
assign CPM[2814] = 12'b111111111111;
assign CPM[2815] = 12'b111111111111;
assign CPM[2816] = 12'b111111111111;
assign CPM[2817] = 12'b111111111111;
assign CPM[2818] = 12'b111111111111;
assign CPM[2819] = 12'b111111111111;
assign CPM[2820] = 12'b000000000000;
assign CPM[2821] = 12'b000000000000;
assign CPM[2822] = 12'b000000000000;
assign CPM[2823] = 12'b000000000000;
assign CPM[2824] = 12'b111111111111;
assign CPM[2825] = 12'b111111111111;
assign CPM[2826] = 12'b111111111111;
assign CPM[2827] = 12'b111111111111;
assign CPM[2828] = 12'b111111111111;
assign CPM[2829] = 12'b111111111111;
assign CPM[2830] = 12'b111111111111;
assign CPM[2831] = 12'b111111111111;
assign CPM[2832] = 12'b111111111111;
assign CPM[2833] = 12'b111111111111;
assign CPM[2834] = 12'b111111111111;
assign CPM[2835] = 12'b111111111111;
assign CPM[2836] = 12'b000000000000;
assign CPM[2837] = 12'b000000000000;
assign CPM[2838] = 12'b000000000000;
assign CPM[2839] = 12'b000000000000;
assign CPM[2840] = 12'b111111111111;
assign CPM[2841] = 12'b111111111111;
assign CPM[2842] = 12'b111111111111;
assign CPM[2843] = 12'b111111111111;
assign CPM[2844] = 12'b111111111111;
assign CPM[2845] = 12'b111111111111;
assign CPM[2846] = 12'b111111111111;
assign CPM[2847] = 12'b111111111111;
assign CPM[2848] = 12'b111111111111;
assign CPM[2849] = 12'b111111111111;
assign CPM[2850] = 12'b111111111111;
assign CPM[2851] = 12'b111111111111;
assign CPM[2852] = 12'b000000000000;
assign CPM[2853] = 12'b000000000000;
assign CPM[2854] = 12'b000000000000;
assign CPM[2855] = 12'b000000000000;
assign CPM[2856] = 12'b111111111111;
assign CPM[2857] = 12'b111111111111;
assign CPM[2858] = 12'b111111111111;
assign CPM[2859] = 12'b111111111111;
assign CPM[2860] = 12'b111111111111;
assign CPM[2861] = 12'b111111111111;
assign CPM[2862] = 12'b111111111111;
assign CPM[2863] = 12'b111111111111;
assign CPM[2864] = 12'b111111111111;
assign CPM[2865] = 12'b111111111111;
assign CPM[2866] = 12'b111111111111;
assign CPM[2867] = 12'b111111111111;
assign CPM[2868] = 12'b000000000000;
assign CPM[2869] = 12'b000000000000;
assign CPM[2870] = 12'b000000000000;
assign CPM[2871] = 12'b000000000000;
assign CPM[2872] = 12'b111111111111;
assign CPM[2873] = 12'b111111111111;
assign CPM[2874] = 12'b111111111111;
assign CPM[2875] = 12'b111111111111;
assign CPM[2876] = 12'b111111111111;
assign CPM[2877] = 12'b111111111111;
assign CPM[2878] = 12'b111111111111;
assign CPM[2879] = 12'b111111111111;
assign CPM[2880] = 12'b111111111111;
assign CPM[2881] = 12'b111111111111;
assign CPM[2882] = 12'b111111111111;
assign CPM[2883] = 12'b111111111111;
assign CPM[2884] = 12'b000000000000;
assign CPM[2885] = 12'b000000000000;
assign CPM[2886] = 12'b000000000000;
assign CPM[2887] = 12'b000000000000;
assign CPM[2888] = 12'b111111111111;
assign CPM[2889] = 12'b111111111111;
assign CPM[2890] = 12'b111111111111;
assign CPM[2891] = 12'b111111111111;
assign CPM[2892] = 12'b111111111111;
assign CPM[2893] = 12'b111111111111;
assign CPM[2894] = 12'b111111111111;
assign CPM[2895] = 12'b111111111111;
assign CPM[2896] = 12'b111111111111;
assign CPM[2897] = 12'b111111111111;
assign CPM[2898] = 12'b111111111111;
assign CPM[2899] = 12'b111111111111;
assign CPM[2900] = 12'b000000000000;
assign CPM[2901] = 12'b000000000000;
assign CPM[2902] = 12'b000000000000;
assign CPM[2903] = 12'b000000000000;
assign CPM[2904] = 12'b111111111111;
assign CPM[2905] = 12'b111111111111;
assign CPM[2906] = 12'b111111111111;
assign CPM[2907] = 12'b111111111111;
assign CPM[2908] = 12'b111111111111;
assign CPM[2909] = 12'b111111111111;
assign CPM[2910] = 12'b111111111111;
assign CPM[2911] = 12'b111111111111;
assign CPM[2912] = 12'b111111111111;
assign CPM[2913] = 12'b111111111111;
assign CPM[2914] = 12'b111111111111;
assign CPM[2915] = 12'b111111111111;
assign CPM[2916] = 12'b000000000000;
assign CPM[2917] = 12'b000000000000;
assign CPM[2918] = 12'b000000000000;
assign CPM[2919] = 12'b000000000000;
assign CPM[2920] = 12'b111111111111;
assign CPM[2921] = 12'b111111111111;
assign CPM[2922] = 12'b111111111111;
assign CPM[2923] = 12'b111111111111;
assign CPM[2924] = 12'b111111111111;
assign CPM[2925] = 12'b111111111111;
assign CPM[2926] = 12'b111111111111;
assign CPM[2927] = 12'b111111111111;
assign CPM[2928] = 12'b111111111111;
assign CPM[2929] = 12'b111111111111;
assign CPM[2930] = 12'b111111111111;
assign CPM[2931] = 12'b111111111111;
assign CPM[2932] = 12'b000000000000;
assign CPM[2933] = 12'b000000000000;
assign CPM[2934] = 12'b000000000000;
assign CPM[2935] = 12'b000000000000;
assign CPM[2936] = 12'b111111111111;
assign CPM[2937] = 12'b111111111111;
assign CPM[2938] = 12'b111111111111;
assign CPM[2939] = 12'b111111111111;
assign CPM[2940] = 12'b111111111111;
assign CPM[2941] = 12'b111111111111;
assign CPM[2942] = 12'b111111111111;
assign CPM[2943] = 12'b111111111111;
assign CPM[2944] = 12'b111111111111;
assign CPM[2945] = 12'b111111111111;
assign CPM[2946] = 12'b111111111111;
assign CPM[2947] = 12'b111111111111;
assign CPM[2948] = 12'b000000000000;
assign CPM[2949] = 12'b000000000000;
assign CPM[2950] = 12'b000000000000;
assign CPM[2951] = 12'b000000000000;
assign CPM[2952] = 12'b111111111111;
assign CPM[2953] = 12'b111111111111;
assign CPM[2954] = 12'b111111111111;
assign CPM[2955] = 12'b111111111111;
assign CPM[2956] = 12'b111111111111;
assign CPM[2957] = 12'b111111111111;
assign CPM[2958] = 12'b111111111111;
assign CPM[2959] = 12'b111111111111;
assign CPM[2960] = 12'b111111111111;
assign CPM[2961] = 12'b111111111111;
assign CPM[2962] = 12'b111111111111;
assign CPM[2963] = 12'b111111111111;
assign CPM[2964] = 12'b000000000000;
assign CPM[2965] = 12'b000000000000;
assign CPM[2966] = 12'b000000000000;
assign CPM[2967] = 12'b000000000000;
assign CPM[2968] = 12'b111111111111;
assign CPM[2969] = 12'b111111111111;
assign CPM[2970] = 12'b111111111111;
assign CPM[2971] = 12'b111111111111;
assign CPM[2972] = 12'b111111111111;
assign CPM[2973] = 12'b111111111111;
assign CPM[2974] = 12'b111111111111;
assign CPM[2975] = 12'b111111111111;
assign CPM[2976] = 12'b111111111111;
assign CPM[2977] = 12'b111111111111;
assign CPM[2978] = 12'b111111111111;
assign CPM[2979] = 12'b111111111111;
assign CPM[2980] = 12'b111111111111;
assign CPM[2981] = 12'b111111111111;
assign CPM[2982] = 12'b111111111111;
assign CPM[2983] = 12'b111111111111;
assign CPM[2984] = 12'b111111111111;
assign CPM[2985] = 12'b111111111111;
assign CPM[2986] = 12'b111111111111;
assign CPM[2987] = 12'b111111111111;
assign CPM[2988] = 12'b111111111111;
assign CPM[2989] = 12'b111111111111;
assign CPM[2990] = 12'b111111111111;
assign CPM[2991] = 12'b111111111111;
assign CPM[2992] = 12'b111111111111;
assign CPM[2993] = 12'b111111111111;
assign CPM[2994] = 12'b111111111111;
assign CPM[2995] = 12'b111111111111;
assign CPM[2996] = 12'b111111111111;
assign CPM[2997] = 12'b111111111111;
assign CPM[2998] = 12'b111111111111;
assign CPM[2999] = 12'b111111111111;
assign CPM[3000] = 12'b111111111111;
assign CPM[3001] = 12'b111111111111;
assign CPM[3002] = 12'b111111111111;
assign CPM[3003] = 12'b111111111111;
assign CPM[3004] = 12'b111111111111;
assign CPM[3005] = 12'b111111111111;
assign CPM[3006] = 12'b111111111111;
assign CPM[3007] = 12'b111111111111;
assign CPM[3008] = 12'b111111111111;
assign CPM[3009] = 12'b111111111111;
assign CPM[3010] = 12'b111111111111;
assign CPM[3011] = 12'b111111111111;
assign CPM[3012] = 12'b111111111111;
assign CPM[3013] = 12'b111111111111;
assign CPM[3014] = 12'b111111111111;
assign CPM[3015] = 12'b111111111111;
assign CPM[3016] = 12'b111111111111;
assign CPM[3017] = 12'b111111111111;
assign CPM[3018] = 12'b111111111111;
assign CPM[3019] = 12'b111111111111;
assign CPM[3020] = 12'b111111111111;
assign CPM[3021] = 12'b111111111111;
assign CPM[3022] = 12'b111111111111;
assign CPM[3023] = 12'b111111111111;
assign CPM[3024] = 12'b111111111111;
assign CPM[3025] = 12'b111111111111;
assign CPM[3026] = 12'b111111111111;
assign CPM[3027] = 12'b111111111111;
assign CPM[3028] = 12'b111111111111;
assign CPM[3029] = 12'b111111111111;
assign CPM[3030] = 12'b111111111111;
assign CPM[3031] = 12'b111111111111;
assign CPM[3032] = 12'b111111111111;
assign CPM[3033] = 12'b111111111111;
assign CPM[3034] = 12'b111111111111;
assign CPM[3035] = 12'b111111111111;
assign CPM[3036] = 12'b111111111111;
assign CPM[3037] = 12'b111111111111;
assign CPM[3038] = 12'b111111111111;
assign CPM[3039] = 12'b111111111111;
assign CPM[3040] = 12'b111111111111;
assign CPM[3041] = 12'b111111111111;
assign CPM[3042] = 12'b111111111111;
assign CPM[3043] = 12'b111111111111;
assign CPM[3044] = 12'b111111111111;
assign CPM[3045] = 12'b111111111111;
assign CPM[3046] = 12'b111111111111;
assign CPM[3047] = 12'b111111111111;
assign CPM[3048] = 12'b111111111111;
assign CPM[3049] = 12'b111111111111;
assign CPM[3050] = 12'b111111111111;
assign CPM[3051] = 12'b111111111111;
assign CPM[3052] = 12'b111111111111;
assign CPM[3053] = 12'b111111111111;
assign CPM[3054] = 12'b111111111111;
assign CPM[3055] = 12'b111111111111;
assign CPM[3056] = 12'b111111111111;
assign CPM[3057] = 12'b111111111111;
assign CPM[3058] = 12'b111111111111;
assign CPM[3059] = 12'b111111111111;
assign CPM[3060] = 12'b111111111111;
assign CPM[3061] = 12'b111111111111;
assign CPM[3062] = 12'b111111111111;
assign CPM[3063] = 12'b111111111111;
assign CPM[3064] = 12'b111111111111;
assign CPM[3065] = 12'b111111111111;
assign CPM[3066] = 12'b111111111111;
assign CPM[3067] = 12'b111111111111;
assign CPM[3068] = 12'b111111111111;
assign CPM[3069] = 12'b111111111111;
assign CPM[3070] = 12'b111111111111;
assign CPM[3071] = 12'b111111111111;
assign CPM[3072] = 12'b111111111111;
assign CPM[3073] = 12'b111111111111;
assign CPM[3074] = 12'b111111111111;
assign CPM[3075] = 12'b111111111111;
assign CPM[3076] = 12'b111111111111;
assign CPM[3077] = 12'b111111111111;
assign CPM[3078] = 12'b111111111111;
assign CPM[3079] = 12'b111111111111;
assign CPM[3080] = 12'b111111111111;
assign CPM[3081] = 12'b111111111111;
assign CPM[3082] = 12'b111111111111;
assign CPM[3083] = 12'b111111111111;
assign CPM[3084] = 12'b111111111111;
assign CPM[3085] = 12'b111111111111;
assign CPM[3086] = 12'b111111111111;
assign CPM[3087] = 12'b111111111111;
assign CPM[3088] = 12'b111111111111;
assign CPM[3089] = 12'b111111111111;
assign CPM[3090] = 12'b111111111111;
assign CPM[3091] = 12'b111111111111;
assign CPM[3092] = 12'b111111111111;
assign CPM[3093] = 12'b111111111111;
assign CPM[3094] = 12'b111111111111;
assign CPM[3095] = 12'b111111111111;
assign CPM[3096] = 12'b111111111111;
assign CPM[3097] = 12'b111111111111;
assign CPM[3098] = 12'b111111111111;
assign CPM[3099] = 12'b111111111111;
assign CPM[3100] = 12'b111111111111;
assign CPM[3101] = 12'b111111111111;
assign CPM[3102] = 12'b111111111111;
assign CPM[3103] = 12'b111111111111;
assign CPM[3104] = 12'b111111111111;
assign CPM[3105] = 12'b111111111111;
assign CPM[3106] = 12'b111111111111;
assign CPM[3107] = 12'b111111111111;
assign CPM[3108] = 12'b111111111111;
assign CPM[3109] = 12'b111111111111;
assign CPM[3110] = 12'b111111111111;
assign CPM[3111] = 12'b111111111111;
assign CPM[3112] = 12'b111111111111;
assign CPM[3113] = 12'b111111111111;
assign CPM[3114] = 12'b111111111111;
assign CPM[3115] = 12'b111111111111;
assign CPM[3116] = 12'b111111111111;
assign CPM[3117] = 12'b111111111111;
assign CPM[3118] = 12'b111111111111;
assign CPM[3119] = 12'b111111111111;
assign CPM[3120] = 12'b111111111111;
assign CPM[3121] = 12'b111111111111;
assign CPM[3122] = 12'b111111111111;
assign CPM[3123] = 12'b111111111111;
assign CPM[3124] = 12'b111111111111;
assign CPM[3125] = 12'b111111111111;
assign CPM[3126] = 12'b111111111111;
assign CPM[3127] = 12'b111111111111;
assign CPM[3128] = 12'b111111111111;
assign CPM[3129] = 12'b111111111111;
assign CPM[3130] = 12'b111111111111;
assign CPM[3131] = 12'b111111111111;
assign CPM[3132] = 12'b111111111111;
assign CPM[3133] = 12'b111111111111;
assign CPM[3134] = 12'b111111111111;
assign CPM[3135] = 12'b111111111111;
assign CPM[3136] = 12'b111111111111;
assign CPM[3137] = 12'b111111111111;
assign CPM[3138] = 12'b111111111111;
assign CPM[3139] = 12'b111111111111;
assign CPM[3140] = 12'b111111111111;
assign CPM[3141] = 12'b111111111111;
assign CPM[3142] = 12'b111111111111;
assign CPM[3143] = 12'b111111111111;
assign CPM[3144] = 12'b111111111111;
assign CPM[3145] = 12'b111111111111;
assign CPM[3146] = 12'b111111111111;
assign CPM[3147] = 12'b111111111111;
assign CPM[3148] = 12'b111111111111;
assign CPM[3149] = 12'b111111111111;
assign CPM[3150] = 12'b111111111111;
assign CPM[3151] = 12'b111111111111;
assign CPM[3152] = 12'b111111111111;
assign CPM[3153] = 12'b111111111111;
assign CPM[3154] = 12'b111111111111;
assign CPM[3155] = 12'b111111111111;
assign CPM[3156] = 12'b111111111111;
assign CPM[3157] = 12'b111111111111;
assign CPM[3158] = 12'b111111111111;
assign CPM[3159] = 12'b111111111111;
assign CPM[3160] = 12'b111111111111;
assign CPM[3161] = 12'b111111111111;
assign CPM[3162] = 12'b111111111111;
assign CPM[3163] = 12'b111111111111;
assign CPM[3164] = 12'b111111111111;
assign CPM[3165] = 12'b111111111111;
assign CPM[3166] = 12'b111111111111;
assign CPM[3167] = 12'b111111111111;
assign CPM[3168] = 12'b111111111111;
assign CPM[3169] = 12'b111111111111;
assign CPM[3170] = 12'b111111111111;
assign CPM[3171] = 12'b111111111111;
assign CPM[3172] = 12'b111111111111;
assign CPM[3173] = 12'b111111111111;
assign CPM[3174] = 12'b111111111111;
assign CPM[3175] = 12'b111111111111;
assign CPM[3176] = 12'b111111111111;
assign CPM[3177] = 12'b000000000000;
assign CPM[3178] = 12'b000000000000;
assign CPM[3179] = 12'b000000000000;
assign CPM[3180] = 12'b000000000000;
assign CPM[3181] = 12'b000000000000;
assign CPM[3182] = 12'b000000000000;
assign CPM[3183] = 12'b000000000000;
assign CPM[3184] = 12'b000000000000;
assign CPM[3185] = 12'b000000000000;
assign CPM[3186] = 12'b000000000000;
assign CPM[3187] = 12'b000000000000;
assign CPM[3188] = 12'b000000000000;
assign CPM[3189] = 12'b000000000000;
assign CPM[3190] = 12'b111111111111;
assign CPM[3191] = 12'b111111111111;
assign CPM[3192] = 12'b111111111111;
assign CPM[3193] = 12'b111111111111;
assign CPM[3194] = 12'b111111111111;
assign CPM[3195] = 12'b111111111111;
assign CPM[3196] = 12'b111111111111;
assign CPM[3197] = 12'b111111111111;
assign CPM[3198] = 12'b111111111111;
assign CPM[3199] = 12'b111111111111;
assign CPM[3200] = 12'b111111111111;
assign CPM[3201] = 12'b111111111111;
assign CPM[3202] = 12'b111111111111;
assign CPM[3203] = 12'b111111111111;
assign CPM[3204] = 12'b111111111111;
assign CPM[3205] = 12'b111111111111;
assign CPM[3206] = 12'b111111111111;
assign CPM[3207] = 12'b111111111111;
assign CPM[3208] = 12'b111111111111;
assign CPM[3209] = 12'b000000000000;
assign CPM[3210] = 12'b000000000000;
assign CPM[3211] = 12'b000000000000;
assign CPM[3212] = 12'b000000000000;
assign CPM[3213] = 12'b000000000000;
assign CPM[3214] = 12'b000000000000;
assign CPM[3215] = 12'b000000000000;
assign CPM[3216] = 12'b000000000000;
assign CPM[3217] = 12'b000000000000;
assign CPM[3218] = 12'b000000000000;
assign CPM[3219] = 12'b000000000000;
assign CPM[3220] = 12'b000000000000;
assign CPM[3221] = 12'b000000000000;
assign CPM[3222] = 12'b111111111111;
assign CPM[3223] = 12'b111111111111;
assign CPM[3224] = 12'b111111111111;
assign CPM[3225] = 12'b111111111111;
assign CPM[3226] = 12'b111111111111;
assign CPM[3227] = 12'b111111111111;
assign CPM[3228] = 12'b111111111111;
assign CPM[3229] = 12'b111111111111;
assign CPM[3230] = 12'b111111111111;
assign CPM[3231] = 12'b111111111111;
assign CPM[3232] = 12'b111111111111;
assign CPM[3233] = 12'b111111111111;
assign CPM[3234] = 12'b111111111111;
assign CPM[3235] = 12'b111111111111;
assign CPM[3236] = 12'b111111111111;
assign CPM[3237] = 12'b111111111111;
assign CPM[3238] = 12'b111111111111;
assign CPM[3239] = 12'b111111111111;
assign CPM[3240] = 12'b111111111111;
assign CPM[3241] = 12'b000000000000;
assign CPM[3242] = 12'b000000000000;
assign CPM[3243] = 12'b000000000000;
assign CPM[3244] = 12'b000000000000;
assign CPM[3245] = 12'b000000000000;
assign CPM[3246] = 12'b000000000000;
assign CPM[3247] = 12'b000000000000;
assign CPM[3248] = 12'b000000000000;
assign CPM[3249] = 12'b000000000000;
assign CPM[3250] = 12'b000000000000;
assign CPM[3251] = 12'b000000000000;
assign CPM[3252] = 12'b000000000000;
assign CPM[3253] = 12'b000000000000;
assign CPM[3254] = 12'b111111111111;
assign CPM[3255] = 12'b111111111111;
assign CPM[3256] = 12'b111111111111;
assign CPM[3257] = 12'b111111111111;
assign CPM[3258] = 12'b111111111111;
assign CPM[3259] = 12'b111111111111;
assign CPM[3260] = 12'b111111111111;
assign CPM[3261] = 12'b111111111111;
assign CPM[3262] = 12'b111111111111;
assign CPM[3263] = 12'b111111111111;
assign CPM[3264] = 12'b111111111111;
assign CPM[3265] = 12'b111111111111;
assign CPM[3266] = 12'b111111111111;
assign CPM[3267] = 12'b111111111111;
assign CPM[3268] = 12'b111111111111;
assign CPM[3269] = 12'b111111111111;
assign CPM[3270] = 12'b111111111111;
assign CPM[3271] = 12'b111111111111;
assign CPM[3272] = 12'b111111111111;
assign CPM[3273] = 12'b000000000000;
assign CPM[3274] = 12'b000000000000;
assign CPM[3275] = 12'b000000000000;
assign CPM[3276] = 12'b000000000000;
assign CPM[3277] = 12'b000000000000;
assign CPM[3278] = 12'b000000000000;
assign CPM[3279] = 12'b000000000000;
assign CPM[3280] = 12'b000000000000;
assign CPM[3281] = 12'b000000000000;
assign CPM[3282] = 12'b000000000000;
assign CPM[3283] = 12'b000000000000;
assign CPM[3284] = 12'b000000000000;
assign CPM[3285] = 12'b000000000000;
assign CPM[3286] = 12'b111111111111;
assign CPM[3287] = 12'b111111111111;
assign CPM[3288] = 12'b111111111111;
assign CPM[3289] = 12'b111111111111;
assign CPM[3290] = 12'b111111111111;
assign CPM[3291] = 12'b111111111111;
assign CPM[3292] = 12'b111111111111;
assign CPM[3293] = 12'b111111111111;
assign CPM[3294] = 12'b111111111111;
assign CPM[3295] = 12'b111111111111;
assign CPM[3296] = 12'b111111111111;
assign CPM[3297] = 12'b111111111111;
assign CPM[3298] = 12'b111111111111;
assign CPM[3299] = 12'b111111111111;
assign CPM[3300] = 12'b111111111111;
assign CPM[3301] = 12'b000000000000;
assign CPM[3302] = 12'b000000000000;
assign CPM[3303] = 12'b000000000000;
assign CPM[3304] = 12'b000000000000;
assign CPM[3305] = 12'b111111111111;
assign CPM[3306] = 12'b111111111111;
assign CPM[3307] = 12'b111111111111;
assign CPM[3308] = 12'b111111111111;
assign CPM[3309] = 12'b111111111111;
assign CPM[3310] = 12'b111111111111;
assign CPM[3311] = 12'b111111111111;
assign CPM[3312] = 12'b111111111111;
assign CPM[3313] = 12'b111111111111;
assign CPM[3314] = 12'b111111111111;
assign CPM[3315] = 12'b111111111111;
assign CPM[3316] = 12'b111111111111;
assign CPM[3317] = 12'b000000000000;
assign CPM[3318] = 12'b000000000000;
assign CPM[3319] = 12'b000000000000;
assign CPM[3320] = 12'b000000000000;
assign CPM[3321] = 12'b111111111111;
assign CPM[3322] = 12'b111111111111;
assign CPM[3323] = 12'b111111111111;
assign CPM[3324] = 12'b111111111111;
assign CPM[3325] = 12'b111111111111;
assign CPM[3326] = 12'b111111111111;
assign CPM[3327] = 12'b111111111111;
assign CPM[3328] = 12'b111111111111;
assign CPM[3329] = 12'b111111111111;
assign CPM[3330] = 12'b111111111111;
assign CPM[3331] = 12'b111111111111;
assign CPM[3332] = 12'b111111111111;
assign CPM[3333] = 12'b000000000000;
assign CPM[3334] = 12'b000000000000;
assign CPM[3335] = 12'b000000000000;
assign CPM[3336] = 12'b000000000000;
assign CPM[3337] = 12'b111111111111;
assign CPM[3338] = 12'b111111111111;
assign CPM[3339] = 12'b111111111111;
assign CPM[3340] = 12'b111111111111;
assign CPM[3341] = 12'b111111111111;
assign CPM[3342] = 12'b111111111111;
assign CPM[3343] = 12'b111111111111;
assign CPM[3344] = 12'b111111111111;
assign CPM[3345] = 12'b111111111111;
assign CPM[3346] = 12'b000000000000;
assign CPM[3347] = 12'b000000000000;
assign CPM[3348] = 12'b000000000000;
assign CPM[3349] = 12'b000000000000;
assign CPM[3350] = 12'b000000000000;
assign CPM[3351] = 12'b000000000000;
assign CPM[3352] = 12'b000000000000;
assign CPM[3353] = 12'b111111111111;
assign CPM[3354] = 12'b111111111111;
assign CPM[3355] = 12'b111111111111;
assign CPM[3356] = 12'b111111111111;
assign CPM[3357] = 12'b111111111111;
assign CPM[3358] = 12'b111111111111;
assign CPM[3359] = 12'b111111111111;
assign CPM[3360] = 12'b111111111111;
assign CPM[3361] = 12'b111111111111;
assign CPM[3362] = 12'b111111111111;
assign CPM[3363] = 12'b111111111111;
assign CPM[3364] = 12'b111111111111;
assign CPM[3365] = 12'b000000000000;
assign CPM[3366] = 12'b000000000000;
assign CPM[3367] = 12'b000000000000;
assign CPM[3368] = 12'b000000000000;
assign CPM[3369] = 12'b111111111111;
assign CPM[3370] = 12'b111111111111;
assign CPM[3371] = 12'b111111111111;
assign CPM[3372] = 12'b111111111111;
assign CPM[3373] = 12'b111111111111;
assign CPM[3374] = 12'b111111111111;
assign CPM[3375] = 12'b111111111111;
assign CPM[3376] = 12'b111111111111;
assign CPM[3377] = 12'b111111111111;
assign CPM[3378] = 12'b000000000000;
assign CPM[3379] = 12'b000000000000;
assign CPM[3380] = 12'b000000000000;
assign CPM[3381] = 12'b000000000000;
assign CPM[3382] = 12'b000000000000;
assign CPM[3383] = 12'b000000000000;
assign CPM[3384] = 12'b000000000000;
assign CPM[3385] = 12'b111111111111;
assign CPM[3386] = 12'b111111111111;
assign CPM[3387] = 12'b111111111111;
assign CPM[3388] = 12'b111111111111;
assign CPM[3389] = 12'b111111111111;
assign CPM[3390] = 12'b111111111111;
assign CPM[3391] = 12'b111111111111;
assign CPM[3392] = 12'b111111111111;
assign CPM[3393] = 12'b111111111111;
assign CPM[3394] = 12'b111111111111;
assign CPM[3395] = 12'b111111111111;
assign CPM[3396] = 12'b111111111111;
assign CPM[3397] = 12'b000000000000;
assign CPM[3398] = 12'b000000000000;
assign CPM[3399] = 12'b000000000000;
assign CPM[3400] = 12'b000000000000;
assign CPM[3401] = 12'b111111111111;
assign CPM[3402] = 12'b111111111111;
assign CPM[3403] = 12'b111111111111;
assign CPM[3404] = 12'b111111111111;
assign CPM[3405] = 12'b111111111111;
assign CPM[3406] = 12'b111111111111;
assign CPM[3407] = 12'b111111111111;
assign CPM[3408] = 12'b111111111111;
assign CPM[3409] = 12'b111111111111;
assign CPM[3410] = 12'b000000000000;
assign CPM[3411] = 12'b000000000000;
assign CPM[3412] = 12'b000000000000;
assign CPM[3413] = 12'b000000000000;
assign CPM[3414] = 12'b000000000000;
assign CPM[3415] = 12'b000000000000;
assign CPM[3416] = 12'b000000000000;
assign CPM[3417] = 12'b111111111111;
assign CPM[3418] = 12'b111111111111;
assign CPM[3419] = 12'b111111111111;
assign CPM[3420] = 12'b111111111111;
assign CPM[3421] = 12'b111111111111;
assign CPM[3422] = 12'b111111111111;
assign CPM[3423] = 12'b111111111111;
assign CPM[3424] = 12'b111111111111;
assign CPM[3425] = 12'b111111111111;
assign CPM[3426] = 12'b111111111111;
assign CPM[3427] = 12'b111111111111;
assign CPM[3428] = 12'b111111111111;
assign CPM[3429] = 12'b000000000000;
assign CPM[3430] = 12'b000000000000;
assign CPM[3431] = 12'b000000000000;
assign CPM[3432] = 12'b000000000000;
assign CPM[3433] = 12'b111111111111;
assign CPM[3434] = 12'b111111111111;
assign CPM[3435] = 12'b111111111111;
assign CPM[3436] = 12'b111111111111;
assign CPM[3437] = 12'b111111111111;
assign CPM[3438] = 12'b111111111111;
assign CPM[3439] = 12'b111111111111;
assign CPM[3440] = 12'b111111111111;
assign CPM[3441] = 12'b111111111111;
assign CPM[3442] = 12'b000000000000;
assign CPM[3443] = 12'b000000000000;
assign CPM[3444] = 12'b000000000000;
assign CPM[3445] = 12'b000000000000;
assign CPM[3446] = 12'b000000000000;
assign CPM[3447] = 12'b000000000000;
assign CPM[3448] = 12'b000000000000;
assign CPM[3449] = 12'b111111111111;
assign CPM[3450] = 12'b111111111111;
assign CPM[3451] = 12'b111111111111;
assign CPM[3452] = 12'b111111111111;
assign CPM[3453] = 12'b111111111111;
assign CPM[3454] = 12'b111111111111;
assign CPM[3455] = 12'b111111111111;
assign CPM[3456] = 12'b111111111111;
assign CPM[3457] = 12'b111111111111;
assign CPM[3458] = 12'b111111111111;
assign CPM[3459] = 12'b111111111111;
assign CPM[3460] = 12'b111111111111;
assign CPM[3461] = 12'b000000000000;
assign CPM[3462] = 12'b000000000000;
assign CPM[3463] = 12'b000000000000;
assign CPM[3464] = 12'b000000000000;
assign CPM[3465] = 12'b111111111111;
assign CPM[3466] = 12'b111111111111;
assign CPM[3467] = 12'b111111111111;
assign CPM[3468] = 12'b111111111111;
assign CPM[3469] = 12'b111111111111;
assign CPM[3470] = 12'b111111111111;
assign CPM[3471] = 12'b000000000000;
assign CPM[3472] = 12'b000000000000;
assign CPM[3473] = 12'b000000000000;
assign CPM[3474] = 12'b111111111111;
assign CPM[3475] = 12'b111111111111;
assign CPM[3476] = 12'b111111111111;
assign CPM[3477] = 12'b000000000000;
assign CPM[3478] = 12'b000000000000;
assign CPM[3479] = 12'b000000000000;
assign CPM[3480] = 12'b000000000000;
assign CPM[3481] = 12'b111111111111;
assign CPM[3482] = 12'b111111111111;
assign CPM[3483] = 12'b111111111111;
assign CPM[3484] = 12'b111111111111;
assign CPM[3485] = 12'b111111111111;
assign CPM[3486] = 12'b111111111111;
assign CPM[3487] = 12'b111111111111;
assign CPM[3488] = 12'b111111111111;
assign CPM[3489] = 12'b111111111111;
assign CPM[3490] = 12'b111111111111;
assign CPM[3491] = 12'b111111111111;
assign CPM[3492] = 12'b111111111111;
assign CPM[3493] = 12'b000000000000;
assign CPM[3494] = 12'b000000000000;
assign CPM[3495] = 12'b000000000000;
assign CPM[3496] = 12'b000000000000;
assign CPM[3497] = 12'b111111111111;
assign CPM[3498] = 12'b111111111111;
assign CPM[3499] = 12'b111111111111;
assign CPM[3500] = 12'b111111111111;
assign CPM[3501] = 12'b111111111111;
assign CPM[3502] = 12'b111111111111;
assign CPM[3503] = 12'b000000000000;
assign CPM[3504] = 12'b000000000000;
assign CPM[3505] = 12'b000000000000;
assign CPM[3506] = 12'b111111111111;
assign CPM[3507] = 12'b111111111111;
assign CPM[3508] = 12'b111111111111;
assign CPM[3509] = 12'b000000000000;
assign CPM[3510] = 12'b000000000000;
assign CPM[3511] = 12'b000000000000;
assign CPM[3512] = 12'b000000000000;
assign CPM[3513] = 12'b111111111111;
assign CPM[3514] = 12'b111111111111;
assign CPM[3515] = 12'b111111111111;
assign CPM[3516] = 12'b111111111111;
assign CPM[3517] = 12'b111111111111;
assign CPM[3518] = 12'b111111111111;
assign CPM[3519] = 12'b111111111111;
assign CPM[3520] = 12'b111111111111;
assign CPM[3521] = 12'b111111111111;
assign CPM[3522] = 12'b111111111111;
assign CPM[3523] = 12'b111111111111;
assign CPM[3524] = 12'b111111111111;
assign CPM[3525] = 12'b000000000000;
assign CPM[3526] = 12'b000000000000;
assign CPM[3527] = 12'b000000000000;
assign CPM[3528] = 12'b000000000000;
assign CPM[3529] = 12'b111111111111;
assign CPM[3530] = 12'b111111111111;
assign CPM[3531] = 12'b111111111111;
assign CPM[3532] = 12'b111111111111;
assign CPM[3533] = 12'b111111111111;
assign CPM[3534] = 12'b111111111111;
assign CPM[3535] = 12'b000000000000;
assign CPM[3536] = 12'b000000000000;
assign CPM[3537] = 12'b000000000000;
assign CPM[3538] = 12'b111111111111;
assign CPM[3539] = 12'b111111111111;
assign CPM[3540] = 12'b111111111111;
assign CPM[3541] = 12'b000000000000;
assign CPM[3542] = 12'b000000000000;
assign CPM[3543] = 12'b000000000000;
assign CPM[3544] = 12'b000000000000;
assign CPM[3545] = 12'b111111111111;
assign CPM[3546] = 12'b111111111111;
assign CPM[3547] = 12'b111111111111;
assign CPM[3548] = 12'b111111111111;
assign CPM[3549] = 12'b111111111111;
assign CPM[3550] = 12'b111111111111;
assign CPM[3551] = 12'b111111111111;
assign CPM[3552] = 12'b111111111111;
assign CPM[3553] = 12'b111111111111;
assign CPM[3554] = 12'b111111111111;
assign CPM[3555] = 12'b111111111111;
assign CPM[3556] = 12'b111111111111;
assign CPM[3557] = 12'b000000000000;
assign CPM[3558] = 12'b000000000000;
assign CPM[3559] = 12'b000000000000;
assign CPM[3560] = 12'b000000000000;
assign CPM[3561] = 12'b111111111111;
assign CPM[3562] = 12'b111111111111;
assign CPM[3563] = 12'b111111111111;
assign CPM[3564] = 12'b111111111111;
assign CPM[3565] = 12'b111111111111;
assign CPM[3566] = 12'b111111111111;
assign CPM[3567] = 12'b000000000000;
assign CPM[3568] = 12'b000000000000;
assign CPM[3569] = 12'b000000000000;
assign CPM[3570] = 12'b111111111111;
assign CPM[3571] = 12'b111111111111;
assign CPM[3572] = 12'b111111111111;
assign CPM[3573] = 12'b000000000000;
assign CPM[3574] = 12'b000000000000;
assign CPM[3575] = 12'b000000000000;
assign CPM[3576] = 12'b000000000000;
assign CPM[3577] = 12'b111111111111;
assign CPM[3578] = 12'b111111111111;
assign CPM[3579] = 12'b111111111111;
assign CPM[3580] = 12'b111111111111;
assign CPM[3581] = 12'b111111111111;
assign CPM[3582] = 12'b111111111111;
assign CPM[3583] = 12'b111111111111;
assign CPM[3584] = 12'b111111111111;
assign CPM[3585] = 12'b111111111111;
assign CPM[3586] = 12'b111111111111;
assign CPM[3587] = 12'b111111111111;
assign CPM[3588] = 12'b111111111111;
assign CPM[3589] = 12'b000000000000;
assign CPM[3590] = 12'b000000000000;
assign CPM[3591] = 12'b000000000000;
assign CPM[3592] = 12'b000000000000;
assign CPM[3593] = 12'b111111111111;
assign CPM[3594] = 12'b111111111111;
assign CPM[3595] = 12'b111111111111;
assign CPM[3596] = 12'b000000000000;
assign CPM[3597] = 12'b000000000000;
assign CPM[3598] = 12'b000000000000;
assign CPM[3599] = 12'b111111111111;
assign CPM[3600] = 12'b111111111111;
assign CPM[3601] = 12'b111111111111;
assign CPM[3602] = 12'b111111111111;
assign CPM[3603] = 12'b111111111111;
assign CPM[3604] = 12'b111111111111;
assign CPM[3605] = 12'b000000000000;
assign CPM[3606] = 12'b000000000000;
assign CPM[3607] = 12'b000000000000;
assign CPM[3608] = 12'b000000000000;
assign CPM[3609] = 12'b111111111111;
assign CPM[3610] = 12'b111111111111;
assign CPM[3611] = 12'b111111111111;
assign CPM[3612] = 12'b111111111111;
assign CPM[3613] = 12'b111111111111;
assign CPM[3614] = 12'b111111111111;
assign CPM[3615] = 12'b111111111111;
assign CPM[3616] = 12'b111111111111;
assign CPM[3617] = 12'b111111111111;
assign CPM[3618] = 12'b111111111111;
assign CPM[3619] = 12'b111111111111;
assign CPM[3620] = 12'b111111111111;
assign CPM[3621] = 12'b000000000000;
assign CPM[3622] = 12'b000000000000;
assign CPM[3623] = 12'b000000000000;
assign CPM[3624] = 12'b000000000000;
assign CPM[3625] = 12'b111111111111;
assign CPM[3626] = 12'b111111111111;
assign CPM[3627] = 12'b111111111111;
assign CPM[3628] = 12'b000000000000;
assign CPM[3629] = 12'b000000000000;
assign CPM[3630] = 12'b000000000000;
assign CPM[3631] = 12'b111111111111;
assign CPM[3632] = 12'b111111111111;
assign CPM[3633] = 12'b111111111111;
assign CPM[3634] = 12'b111111111111;
assign CPM[3635] = 12'b111111111111;
assign CPM[3636] = 12'b111111111111;
assign CPM[3637] = 12'b000000000000;
assign CPM[3638] = 12'b000000000000;
assign CPM[3639] = 12'b000000000000;
assign CPM[3640] = 12'b000000000000;
assign CPM[3641] = 12'b111111111111;
assign CPM[3642] = 12'b111111111111;
assign CPM[3643] = 12'b111111111111;
assign CPM[3644] = 12'b111111111111;
assign CPM[3645] = 12'b111111111111;
assign CPM[3646] = 12'b111111111111;
assign CPM[3647] = 12'b111111111111;
assign CPM[3648] = 12'b111111111111;
assign CPM[3649] = 12'b111111111111;
assign CPM[3650] = 12'b111111111111;
assign CPM[3651] = 12'b111111111111;
assign CPM[3652] = 12'b111111111111;
assign CPM[3653] = 12'b000000000000;
assign CPM[3654] = 12'b000000000000;
assign CPM[3655] = 12'b000000000000;
assign CPM[3656] = 12'b000000000000;
assign CPM[3657] = 12'b111111111111;
assign CPM[3658] = 12'b111111111111;
assign CPM[3659] = 12'b111111111111;
assign CPM[3660] = 12'b000000000000;
assign CPM[3661] = 12'b000000000000;
assign CPM[3662] = 12'b000000000000;
assign CPM[3663] = 12'b111111111111;
assign CPM[3664] = 12'b111111111111;
assign CPM[3665] = 12'b111111111111;
assign CPM[3666] = 12'b111111111111;
assign CPM[3667] = 12'b111111111111;
assign CPM[3668] = 12'b111111111111;
assign CPM[3669] = 12'b000000000000;
assign CPM[3670] = 12'b000000000000;
assign CPM[3671] = 12'b000000000000;
assign CPM[3672] = 12'b000000000000;
assign CPM[3673] = 12'b111111111111;
assign CPM[3674] = 12'b111111111111;
assign CPM[3675] = 12'b111111111111;
assign CPM[3676] = 12'b111111111111;
assign CPM[3677] = 12'b111111111111;
assign CPM[3678] = 12'b111111111111;
assign CPM[3679] = 12'b111111111111;
assign CPM[3680] = 12'b111111111111;
assign CPM[3681] = 12'b111111111111;
assign CPM[3682] = 12'b111111111111;
assign CPM[3683] = 12'b111111111111;
assign CPM[3684] = 12'b111111111111;
assign CPM[3685] = 12'b000000000000;
assign CPM[3686] = 12'b000000000000;
assign CPM[3687] = 12'b000000000000;
assign CPM[3688] = 12'b000000000000;
assign CPM[3689] = 12'b111111111111;
assign CPM[3690] = 12'b111111111111;
assign CPM[3691] = 12'b111111111111;
assign CPM[3692] = 12'b000000000000;
assign CPM[3693] = 12'b000000000000;
assign CPM[3694] = 12'b000000000000;
assign CPM[3695] = 12'b111111111111;
assign CPM[3696] = 12'b111111111111;
assign CPM[3697] = 12'b111111111111;
assign CPM[3698] = 12'b111111111111;
assign CPM[3699] = 12'b111111111111;
assign CPM[3700] = 12'b111111111111;
assign CPM[3701] = 12'b000000000000;
assign CPM[3702] = 12'b000000000000;
assign CPM[3703] = 12'b000000000000;
assign CPM[3704] = 12'b000000000000;
assign CPM[3705] = 12'b111111111111;
assign CPM[3706] = 12'b111111111111;
assign CPM[3707] = 12'b111111111111;
assign CPM[3708] = 12'b111111111111;
assign CPM[3709] = 12'b111111111111;
assign CPM[3710] = 12'b111111111111;
assign CPM[3711] = 12'b111111111111;
assign CPM[3712] = 12'b111111111111;
assign CPM[3713] = 12'b111111111111;
assign CPM[3714] = 12'b111111111111;
assign CPM[3715] = 12'b111111111111;
assign CPM[3716] = 12'b111111111111;
assign CPM[3717] = 12'b000000000000;
assign CPM[3718] = 12'b000000000000;
assign CPM[3719] = 12'b000000000000;
assign CPM[3720] = 12'b000000000000;
assign CPM[3721] = 12'b000000000000;
assign CPM[3722] = 12'b000000000000;
assign CPM[3723] = 12'b000000000000;
assign CPM[3724] = 12'b111111111111;
assign CPM[3725] = 12'b111111111111;
assign CPM[3726] = 12'b111111111111;
assign CPM[3727] = 12'b111111111111;
assign CPM[3728] = 12'b111111111111;
assign CPM[3729] = 12'b111111111111;
assign CPM[3730] = 12'b111111111111;
assign CPM[3731] = 12'b111111111111;
assign CPM[3732] = 12'b111111111111;
assign CPM[3733] = 12'b000000000000;
assign CPM[3734] = 12'b000000000000;
assign CPM[3735] = 12'b000000000000;
assign CPM[3736] = 12'b000000000000;
assign CPM[3737] = 12'b111111111111;
assign CPM[3738] = 12'b111111111111;
assign CPM[3739] = 12'b111111111111;
assign CPM[3740] = 12'b111111111111;
assign CPM[3741] = 12'b111111111111;
assign CPM[3742] = 12'b111111111111;
assign CPM[3743] = 12'b111111111111;
assign CPM[3744] = 12'b111111111111;
assign CPM[3745] = 12'b111111111111;
assign CPM[3746] = 12'b111111111111;
assign CPM[3747] = 12'b111111111111;
assign CPM[3748] = 12'b111111111111;
assign CPM[3749] = 12'b000000000000;
assign CPM[3750] = 12'b000000000000;
assign CPM[3751] = 12'b000000000000;
assign CPM[3752] = 12'b000000000000;
assign CPM[3753] = 12'b000000000000;
assign CPM[3754] = 12'b000000000000;
assign CPM[3755] = 12'b000000000000;
assign CPM[3756] = 12'b111111111111;
assign CPM[3757] = 12'b111111111111;
assign CPM[3758] = 12'b111111111111;
assign CPM[3759] = 12'b111111111111;
assign CPM[3760] = 12'b111111111111;
assign CPM[3761] = 12'b111111111111;
assign CPM[3762] = 12'b111111111111;
assign CPM[3763] = 12'b111111111111;
assign CPM[3764] = 12'b111111111111;
assign CPM[3765] = 12'b000000000000;
assign CPM[3766] = 12'b000000000000;
assign CPM[3767] = 12'b000000000000;
assign CPM[3768] = 12'b000000000000;
assign CPM[3769] = 12'b111111111111;
assign CPM[3770] = 12'b111111111111;
assign CPM[3771] = 12'b111111111111;
assign CPM[3772] = 12'b111111111111;
assign CPM[3773] = 12'b111111111111;
assign CPM[3774] = 12'b111111111111;
assign CPM[3775] = 12'b111111111111;
assign CPM[3776] = 12'b111111111111;
assign CPM[3777] = 12'b111111111111;
assign CPM[3778] = 12'b111111111111;
assign CPM[3779] = 12'b111111111111;
assign CPM[3780] = 12'b111111111111;
assign CPM[3781] = 12'b000000000000;
assign CPM[3782] = 12'b000000000000;
assign CPM[3783] = 12'b000000000000;
assign CPM[3784] = 12'b000000000000;
assign CPM[3785] = 12'b000000000000;
assign CPM[3786] = 12'b000000000000;
assign CPM[3787] = 12'b000000000000;
assign CPM[3788] = 12'b111111111111;
assign CPM[3789] = 12'b111111111111;
assign CPM[3790] = 12'b111111111111;
assign CPM[3791] = 12'b111111111111;
assign CPM[3792] = 12'b111111111111;
assign CPM[3793] = 12'b111111111111;
assign CPM[3794] = 12'b111111111111;
assign CPM[3795] = 12'b111111111111;
assign CPM[3796] = 12'b111111111111;
assign CPM[3797] = 12'b000000000000;
assign CPM[3798] = 12'b000000000000;
assign CPM[3799] = 12'b000000000000;
assign CPM[3800] = 12'b000000000000;
assign CPM[3801] = 12'b111111111111;
assign CPM[3802] = 12'b111111111111;
assign CPM[3803] = 12'b111111111111;
assign CPM[3804] = 12'b111111111111;
assign CPM[3805] = 12'b111111111111;
assign CPM[3806] = 12'b111111111111;
assign CPM[3807] = 12'b111111111111;
assign CPM[3808] = 12'b111111111111;
assign CPM[3809] = 12'b111111111111;
assign CPM[3810] = 12'b111111111111;
assign CPM[3811] = 12'b111111111111;
assign CPM[3812] = 12'b111111111111;
assign CPM[3813] = 12'b000000000000;
assign CPM[3814] = 12'b000000000000;
assign CPM[3815] = 12'b000000000000;
assign CPM[3816] = 12'b000000000000;
assign CPM[3817] = 12'b000000000000;
assign CPM[3818] = 12'b000000000000;
assign CPM[3819] = 12'b000000000000;
assign CPM[3820] = 12'b111111111111;
assign CPM[3821] = 12'b111111111111;
assign CPM[3822] = 12'b111111111111;
assign CPM[3823] = 12'b111111111111;
assign CPM[3824] = 12'b111111111111;
assign CPM[3825] = 12'b111111111111;
assign CPM[3826] = 12'b111111111111;
assign CPM[3827] = 12'b111111111111;
assign CPM[3828] = 12'b111111111111;
assign CPM[3829] = 12'b000000000000;
assign CPM[3830] = 12'b000000000000;
assign CPM[3831] = 12'b000000000000;
assign CPM[3832] = 12'b000000000000;
assign CPM[3833] = 12'b111111111111;
assign CPM[3834] = 12'b111111111111;
assign CPM[3835] = 12'b111111111111;
assign CPM[3836] = 12'b111111111111;
assign CPM[3837] = 12'b111111111111;
assign CPM[3838] = 12'b111111111111;
assign CPM[3839] = 12'b111111111111;
assign CPM[3840] = 12'b111111111111;
assign CPM[3841] = 12'b111111111111;
assign CPM[3842] = 12'b111111111111;
assign CPM[3843] = 12'b111111111111;
assign CPM[3844] = 12'b111111111111;
assign CPM[3845] = 12'b000000000000;
assign CPM[3846] = 12'b000000000000;
assign CPM[3847] = 12'b000000000000;
assign CPM[3848] = 12'b000000000000;
assign CPM[3849] = 12'b111111111111;
assign CPM[3850] = 12'b111111111111;
assign CPM[3851] = 12'b111111111111;
assign CPM[3852] = 12'b111111111111;
assign CPM[3853] = 12'b111111111111;
assign CPM[3854] = 12'b111111111111;
assign CPM[3855] = 12'b111111111111;
assign CPM[3856] = 12'b111111111111;
assign CPM[3857] = 12'b111111111111;
assign CPM[3858] = 12'b111111111111;
assign CPM[3859] = 12'b111111111111;
assign CPM[3860] = 12'b111111111111;
assign CPM[3861] = 12'b000000000000;
assign CPM[3862] = 12'b000000000000;
assign CPM[3863] = 12'b000000000000;
assign CPM[3864] = 12'b000000000000;
assign CPM[3865] = 12'b111111111111;
assign CPM[3866] = 12'b111111111111;
assign CPM[3867] = 12'b111111111111;
assign CPM[3868] = 12'b111111111111;
assign CPM[3869] = 12'b111111111111;
assign CPM[3870] = 12'b111111111111;
assign CPM[3871] = 12'b111111111111;
assign CPM[3872] = 12'b111111111111;
assign CPM[3873] = 12'b111111111111;
assign CPM[3874] = 12'b111111111111;
assign CPM[3875] = 12'b111111111111;
assign CPM[3876] = 12'b111111111111;
assign CPM[3877] = 12'b000000000000;
assign CPM[3878] = 12'b000000000000;
assign CPM[3879] = 12'b000000000000;
assign CPM[3880] = 12'b000000000000;
assign CPM[3881] = 12'b111111111111;
assign CPM[3882] = 12'b111111111111;
assign CPM[3883] = 12'b111111111111;
assign CPM[3884] = 12'b111111111111;
assign CPM[3885] = 12'b111111111111;
assign CPM[3886] = 12'b111111111111;
assign CPM[3887] = 12'b111111111111;
assign CPM[3888] = 12'b111111111111;
assign CPM[3889] = 12'b111111111111;
assign CPM[3890] = 12'b111111111111;
assign CPM[3891] = 12'b111111111111;
assign CPM[3892] = 12'b111111111111;
assign CPM[3893] = 12'b000000000000;
assign CPM[3894] = 12'b000000000000;
assign CPM[3895] = 12'b000000000000;
assign CPM[3896] = 12'b000000000000;
assign CPM[3897] = 12'b111111111111;
assign CPM[3898] = 12'b111111111111;
assign CPM[3899] = 12'b111111111111;
assign CPM[3900] = 12'b111111111111;
assign CPM[3901] = 12'b111111111111;
assign CPM[3902] = 12'b111111111111;
assign CPM[3903] = 12'b111111111111;
assign CPM[3904] = 12'b111111111111;
assign CPM[3905] = 12'b111111111111;
assign CPM[3906] = 12'b111111111111;
assign CPM[3907] = 12'b111111111111;
assign CPM[3908] = 12'b111111111111;
assign CPM[3909] = 12'b111111111111;
assign CPM[3910] = 12'b111111111111;
assign CPM[3911] = 12'b111111111111;
assign CPM[3912] = 12'b111111111111;
assign CPM[3913] = 12'b000000000000;
assign CPM[3914] = 12'b000000000000;
assign CPM[3915] = 12'b000000000000;
assign CPM[3916] = 12'b000000000000;
assign CPM[3917] = 12'b000000000000;
assign CPM[3918] = 12'b000000000000;
assign CPM[3919] = 12'b000000000000;
assign CPM[3920] = 12'b000000000000;
assign CPM[3921] = 12'b000000000000;
assign CPM[3922] = 12'b000000000000;
assign CPM[3923] = 12'b000000000000;
assign CPM[3924] = 12'b000000000000;
assign CPM[3925] = 12'b000000000000;
assign CPM[3926] = 12'b111111111111;
assign CPM[3927] = 12'b111111111111;
assign CPM[3928] = 12'b111111111111;
assign CPM[3929] = 12'b111111111111;
assign CPM[3930] = 12'b111111111111;
assign CPM[3931] = 12'b111111111111;
assign CPM[3932] = 12'b111111111111;
assign CPM[3933] = 12'b111111111111;
assign CPM[3934] = 12'b111111111111;
assign CPM[3935] = 12'b111111111111;
assign CPM[3936] = 12'b111111111111;
assign CPM[3937] = 12'b111111111111;
assign CPM[3938] = 12'b111111111111;
assign CPM[3939] = 12'b111111111111;
assign CPM[3940] = 12'b111111111111;
assign CPM[3941] = 12'b111111111111;
assign CPM[3942] = 12'b111111111111;
assign CPM[3943] = 12'b111111111111;
assign CPM[3944] = 12'b111111111111;
assign CPM[3945] = 12'b000000000000;
assign CPM[3946] = 12'b000000000000;
assign CPM[3947] = 12'b000000000000;
assign CPM[3948] = 12'b000000000000;
assign CPM[3949] = 12'b000000000000;
assign CPM[3950] = 12'b000000000000;
assign CPM[3951] = 12'b000000000000;
assign CPM[3952] = 12'b000000000000;
assign CPM[3953] = 12'b000000000000;
assign CPM[3954] = 12'b000000000000;
assign CPM[3955] = 12'b000000000000;
assign CPM[3956] = 12'b000000000000;
assign CPM[3957] = 12'b000000000000;
assign CPM[3958] = 12'b111111111111;
assign CPM[3959] = 12'b111111111111;
assign CPM[3960] = 12'b111111111111;
assign CPM[3961] = 12'b111111111111;
assign CPM[3962] = 12'b111111111111;
assign CPM[3963] = 12'b111111111111;
assign CPM[3964] = 12'b111111111111;
assign CPM[3965] = 12'b111111111111;
assign CPM[3966] = 12'b111111111111;
assign CPM[3967] = 12'b111111111111;
assign CPM[3968] = 12'b111111111111;
assign CPM[3969] = 12'b111111111111;
assign CPM[3970] = 12'b111111111111;
assign CPM[3971] = 12'b111111111111;
assign CPM[3972] = 12'b111111111111;
assign CPM[3973] = 12'b111111111111;
assign CPM[3974] = 12'b111111111111;
assign CPM[3975] = 12'b111111111111;
assign CPM[3976] = 12'b111111111111;
assign CPM[3977] = 12'b000000000000;
assign CPM[3978] = 12'b000000000000;
assign CPM[3979] = 12'b000000000000;
assign CPM[3980] = 12'b000000000000;
assign CPM[3981] = 12'b000000000000;
assign CPM[3982] = 12'b000000000000;
assign CPM[3983] = 12'b000000000000;
assign CPM[3984] = 12'b000000000000;
assign CPM[3985] = 12'b000000000000;
assign CPM[3986] = 12'b000000000000;
assign CPM[3987] = 12'b000000000000;
assign CPM[3988] = 12'b000000000000;
assign CPM[3989] = 12'b000000000000;
assign CPM[3990] = 12'b111111111111;
assign CPM[3991] = 12'b111111111111;
assign CPM[3992] = 12'b111111111111;
assign CPM[3993] = 12'b111111111111;
assign CPM[3994] = 12'b111111111111;
assign CPM[3995] = 12'b111111111111;
assign CPM[3996] = 12'b111111111111;
assign CPM[3997] = 12'b111111111111;
assign CPM[3998] = 12'b111111111111;
assign CPM[3999] = 12'b111111111111;
assign CPM[4000] = 12'b111111111111;
assign CPM[4001] = 12'b111111111111;
assign CPM[4002] = 12'b111111111111;
assign CPM[4003] = 12'b111111111111;
assign CPM[4004] = 12'b111111111111;
assign CPM[4005] = 12'b111111111111;
assign CPM[4006] = 12'b111111111111;
assign CPM[4007] = 12'b111111111111;
assign CPM[4008] = 12'b111111111111;
assign CPM[4009] = 12'b000000000000;
assign CPM[4010] = 12'b000000000000;
assign CPM[4011] = 12'b000000000000;
assign CPM[4012] = 12'b000000000000;
assign CPM[4013] = 12'b000000000000;
assign CPM[4014] = 12'b000000000000;
assign CPM[4015] = 12'b000000000000;
assign CPM[4016] = 12'b000000000000;
assign CPM[4017] = 12'b000000000000;
assign CPM[4018] = 12'b000000000000;
assign CPM[4019] = 12'b000000000000;
assign CPM[4020] = 12'b000000000000;
assign CPM[4021] = 12'b000000000000;
assign CPM[4022] = 12'b111111111111;
assign CPM[4023] = 12'b111111111111;
assign CPM[4024] = 12'b111111111111;
assign CPM[4025] = 12'b111111111111;
assign CPM[4026] = 12'b111111111111;
assign CPM[4027] = 12'b111111111111;
assign CPM[4028] = 12'b111111111111;
assign CPM[4029] = 12'b111111111111;
assign CPM[4030] = 12'b111111111111;
assign CPM[4031] = 12'b111111111111;
assign CPM[4032] = 12'b111111111111;
assign CPM[4033] = 12'b111111111111;
assign CPM[4034] = 12'b111111111111;
assign CPM[4035] = 12'b111111111111;
assign CPM[4036] = 12'b111111111111;
assign CPM[4037] = 12'b111111111111;
assign CPM[4038] = 12'b111111111111;
assign CPM[4039] = 12'b111111111111;
assign CPM[4040] = 12'b111111111111;
assign CPM[4041] = 12'b111111111111;
assign CPM[4042] = 12'b111111111111;
assign CPM[4043] = 12'b111111111111;
assign CPM[4044] = 12'b111111111111;
assign CPM[4045] = 12'b111111111111;
assign CPM[4046] = 12'b111111111111;
assign CPM[4047] = 12'b111111111111;
assign CPM[4048] = 12'b111111111111;
assign CPM[4049] = 12'b111111111111;
assign CPM[4050] = 12'b111111111111;
assign CPM[4051] = 12'b111111111111;
assign CPM[4052] = 12'b111111111111;
assign CPM[4053] = 12'b111111111111;
assign CPM[4054] = 12'b111111111111;
assign CPM[4055] = 12'b111111111111;
assign CPM[4056] = 12'b111111111111;
assign CPM[4057] = 12'b111111111111;
assign CPM[4058] = 12'b111111111111;
assign CPM[4059] = 12'b111111111111;
assign CPM[4060] = 12'b111111111111;
assign CPM[4061] = 12'b111111111111;
assign CPM[4062] = 12'b111111111111;
assign CPM[4063] = 12'b111111111111;
assign CPM[4064] = 12'b111111111111;
assign CPM[4065] = 12'b111111111111;
assign CPM[4066] = 12'b111111111111;
assign CPM[4067] = 12'b111111111111;
assign CPM[4068] = 12'b111111111111;
assign CPM[4069] = 12'b111111111111;
assign CPM[4070] = 12'b111111111111;
assign CPM[4071] = 12'b111111111111;
assign CPM[4072] = 12'b111111111111;
assign CPM[4073] = 12'b111111111111;
assign CPM[4074] = 12'b111111111111;
assign CPM[4075] = 12'b111111111111;
assign CPM[4076] = 12'b111111111111;
assign CPM[4077] = 12'b111111111111;
assign CPM[4078] = 12'b111111111111;
assign CPM[4079] = 12'b111111111111;
assign CPM[4080] = 12'b111111111111;
assign CPM[4081] = 12'b111111111111;
assign CPM[4082] = 12'b111111111111;
assign CPM[4083] = 12'b111111111111;
assign CPM[4084] = 12'b111111111111;
assign CPM[4085] = 12'b111111111111;
assign CPM[4086] = 12'b111111111111;
assign CPM[4087] = 12'b111111111111;
assign CPM[4088] = 12'b111111111111;
assign CPM[4089] = 12'b111111111111;
assign CPM[4090] = 12'b111111111111;
assign CPM[4091] = 12'b111111111111;
assign CPM[4092] = 12'b111111111111;
assign CPM[4093] = 12'b111111111111;
assign CPM[4094] = 12'b111111111111;
assign CPM[4095] = 12'b111111111111;
assign CPM[4096] = 12'b111111111111;
assign CPM[4097] = 12'b111111111111;
assign CPM[4098] = 12'b111111111111;
assign CPM[4099] = 12'b111111111111;
assign CPM[4100] = 12'b111111111111;
assign CPM[4101] = 12'b111111111111;
assign CPM[4102] = 12'b111111111111;
assign CPM[4103] = 12'b111111111111;
assign CPM[4104] = 12'b111111111111;
assign CPM[4105] = 12'b111111111111;
assign CPM[4106] = 12'b111111111111;
assign CPM[4107] = 12'b111111111111;
assign CPM[4108] = 12'b111111111111;
assign CPM[4109] = 12'b111111111111;
assign CPM[4110] = 12'b111111111111;
assign CPM[4111] = 12'b111111111111;
assign CPM[4112] = 12'b111111111111;
assign CPM[4113] = 12'b111111111111;
assign CPM[4114] = 12'b111111111111;
assign CPM[4115] = 12'b111111111111;
assign CPM[4116] = 12'b111111111111;
assign CPM[4117] = 12'b111111111111;
assign CPM[4118] = 12'b111111111111;
assign CPM[4119] = 12'b111111111111;
assign CPM[4120] = 12'b111111111111;
assign CPM[4121] = 12'b111111111111;
assign CPM[4122] = 12'b111111111111;
assign CPM[4123] = 12'b111111111111;
assign CPM[4124] = 12'b111111111111;
assign CPM[4125] = 12'b111111111111;
assign CPM[4126] = 12'b111111111111;
assign CPM[4127] = 12'b111111111111;
assign CPM[4128] = 12'b111111111111;
assign CPM[4129] = 12'b111111111111;
assign CPM[4130] = 12'b111111111111;
assign CPM[4131] = 12'b111111111111;
assign CPM[4132] = 12'b111111111111;
assign CPM[4133] = 12'b111111111111;
assign CPM[4134] = 12'b111111111111;
assign CPM[4135] = 12'b111111111111;
assign CPM[4136] = 12'b111111111111;
assign CPM[4137] = 12'b111111111111;
assign CPM[4138] = 12'b111111111111;
assign CPM[4139] = 12'b111111111111;
assign CPM[4140] = 12'b111111111111;
assign CPM[4141] = 12'b111111111111;
assign CPM[4142] = 12'b111111111111;
assign CPM[4143] = 12'b111111111111;
assign CPM[4144] = 12'b111111111111;
assign CPM[4145] = 12'b111111111111;
assign CPM[4146] = 12'b111111111111;
assign CPM[4147] = 12'b111111111111;
assign CPM[4148] = 12'b111111111111;
assign CPM[4149] = 12'b111111111111;
assign CPM[4150] = 12'b111111111111;
assign CPM[4151] = 12'b111111111111;
assign CPM[4152] = 12'b111111111111;
assign CPM[4153] = 12'b111111111111;
assign CPM[4154] = 12'b111111111111;
assign CPM[4155] = 12'b111111111111;
assign CPM[4156] = 12'b111111111111;
assign CPM[4157] = 12'b111111111111;
assign CPM[4158] = 12'b111111111111;
assign CPM[4159] = 12'b111111111111;
assign CPM[4160] = 12'b111111111111;
assign CPM[4161] = 12'b111111111111;
assign CPM[4162] = 12'b111111111111;
assign CPM[4163] = 12'b111111111111;
assign CPM[4164] = 12'b111111111111;
assign CPM[4165] = 12'b111111111111;
assign CPM[4166] = 12'b111111111111;
assign CPM[4167] = 12'b111111111111;
assign CPM[4168] = 12'b111111111111;
assign CPM[4169] = 12'b111111111111;
assign CPM[4170] = 12'b111111111111;
assign CPM[4171] = 12'b111111111111;
assign CPM[4172] = 12'b111111111111;
assign CPM[4173] = 12'b111111111111;
assign CPM[4174] = 12'b111111111111;
assign CPM[4175] = 12'b000000000000;
assign CPM[4176] = 12'b000000000000;
assign CPM[4177] = 12'b000000000000;
assign CPM[4178] = 12'b000000000000;
assign CPM[4179] = 12'b111111111111;
assign CPM[4180] = 12'b111111111111;
assign CPM[4181] = 12'b111111111111;
assign CPM[4182] = 12'b111111111111;
assign CPM[4183] = 12'b111111111111;
assign CPM[4184] = 12'b111111111111;
assign CPM[4185] = 12'b111111111111;
assign CPM[4186] = 12'b111111111111;
assign CPM[4187] = 12'b111111111111;
assign CPM[4188] = 12'b111111111111;
assign CPM[4189] = 12'b111111111111;
assign CPM[4190] = 12'b111111111111;
assign CPM[4191] = 12'b111111111111;
assign CPM[4192] = 12'b111111111111;
assign CPM[4193] = 12'b111111111111;
assign CPM[4194] = 12'b111111111111;
assign CPM[4195] = 12'b111111111111;
assign CPM[4196] = 12'b111111111111;
assign CPM[4197] = 12'b111111111111;
assign CPM[4198] = 12'b111111111111;
assign CPM[4199] = 12'b111111111111;
assign CPM[4200] = 12'b111111111111;
assign CPM[4201] = 12'b111111111111;
assign CPM[4202] = 12'b111111111111;
assign CPM[4203] = 12'b111111111111;
assign CPM[4204] = 12'b111111111111;
assign CPM[4205] = 12'b111111111111;
assign CPM[4206] = 12'b111111111111;
assign CPM[4207] = 12'b000000000000;
assign CPM[4208] = 12'b000000000000;
assign CPM[4209] = 12'b000000000000;
assign CPM[4210] = 12'b000000000000;
assign CPM[4211] = 12'b111111111111;
assign CPM[4212] = 12'b111111111111;
assign CPM[4213] = 12'b111111111111;
assign CPM[4214] = 12'b111111111111;
assign CPM[4215] = 12'b111111111111;
assign CPM[4216] = 12'b111111111111;
assign CPM[4217] = 12'b111111111111;
assign CPM[4218] = 12'b111111111111;
assign CPM[4219] = 12'b111111111111;
assign CPM[4220] = 12'b111111111111;
assign CPM[4221] = 12'b111111111111;
assign CPM[4222] = 12'b111111111111;
assign CPM[4223] = 12'b111111111111;
assign CPM[4224] = 12'b111111111111;
assign CPM[4225] = 12'b111111111111;
assign CPM[4226] = 12'b111111111111;
assign CPM[4227] = 12'b111111111111;
assign CPM[4228] = 12'b111111111111;
assign CPM[4229] = 12'b111111111111;
assign CPM[4230] = 12'b111111111111;
assign CPM[4231] = 12'b111111111111;
assign CPM[4232] = 12'b111111111111;
assign CPM[4233] = 12'b111111111111;
assign CPM[4234] = 12'b111111111111;
assign CPM[4235] = 12'b111111111111;
assign CPM[4236] = 12'b111111111111;
assign CPM[4237] = 12'b111111111111;
assign CPM[4238] = 12'b111111111111;
assign CPM[4239] = 12'b000000000000;
assign CPM[4240] = 12'b000000000000;
assign CPM[4241] = 12'b000000000000;
assign CPM[4242] = 12'b000000000000;
assign CPM[4243] = 12'b111111111111;
assign CPM[4244] = 12'b111111111111;
assign CPM[4245] = 12'b111111111111;
assign CPM[4246] = 12'b111111111111;
assign CPM[4247] = 12'b111111111111;
assign CPM[4248] = 12'b111111111111;
assign CPM[4249] = 12'b111111111111;
assign CPM[4250] = 12'b111111111111;
assign CPM[4251] = 12'b111111111111;
assign CPM[4252] = 12'b111111111111;
assign CPM[4253] = 12'b111111111111;
assign CPM[4254] = 12'b111111111111;
assign CPM[4255] = 12'b111111111111;
assign CPM[4256] = 12'b111111111111;
assign CPM[4257] = 12'b111111111111;
assign CPM[4258] = 12'b111111111111;
assign CPM[4259] = 12'b111111111111;
assign CPM[4260] = 12'b111111111111;
assign CPM[4261] = 12'b111111111111;
assign CPM[4262] = 12'b111111111111;
assign CPM[4263] = 12'b111111111111;
assign CPM[4264] = 12'b111111111111;
assign CPM[4265] = 12'b111111111111;
assign CPM[4266] = 12'b111111111111;
assign CPM[4267] = 12'b000000000000;
assign CPM[4268] = 12'b000000000000;
assign CPM[4269] = 12'b000000000000;
assign CPM[4270] = 12'b000000000000;
assign CPM[4271] = 12'b000000000000;
assign CPM[4272] = 12'b000000000000;
assign CPM[4273] = 12'b000000000000;
assign CPM[4274] = 12'b000000000000;
assign CPM[4275] = 12'b111111111111;
assign CPM[4276] = 12'b111111111111;
assign CPM[4277] = 12'b111111111111;
assign CPM[4278] = 12'b111111111111;
assign CPM[4279] = 12'b111111111111;
assign CPM[4280] = 12'b111111111111;
assign CPM[4281] = 12'b111111111111;
assign CPM[4282] = 12'b111111111111;
assign CPM[4283] = 12'b111111111111;
assign CPM[4284] = 12'b111111111111;
assign CPM[4285] = 12'b111111111111;
assign CPM[4286] = 12'b111111111111;
assign CPM[4287] = 12'b111111111111;
assign CPM[4288] = 12'b111111111111;
assign CPM[4289] = 12'b111111111111;
assign CPM[4290] = 12'b111111111111;
assign CPM[4291] = 12'b111111111111;
assign CPM[4292] = 12'b111111111111;
assign CPM[4293] = 12'b111111111111;
assign CPM[4294] = 12'b111111111111;
assign CPM[4295] = 12'b111111111111;
assign CPM[4296] = 12'b111111111111;
assign CPM[4297] = 12'b111111111111;
assign CPM[4298] = 12'b111111111111;
assign CPM[4299] = 12'b000000000000;
assign CPM[4300] = 12'b000000000000;
assign CPM[4301] = 12'b000000000000;
assign CPM[4302] = 12'b000000000000;
assign CPM[4303] = 12'b000000000000;
assign CPM[4304] = 12'b000000000000;
assign CPM[4305] = 12'b000000000000;
assign CPM[4306] = 12'b000000000000;
assign CPM[4307] = 12'b111111111111;
assign CPM[4308] = 12'b111111111111;
assign CPM[4309] = 12'b111111111111;
assign CPM[4310] = 12'b111111111111;
assign CPM[4311] = 12'b111111111111;
assign CPM[4312] = 12'b111111111111;
assign CPM[4313] = 12'b111111111111;
assign CPM[4314] = 12'b111111111111;
assign CPM[4315] = 12'b111111111111;
assign CPM[4316] = 12'b111111111111;
assign CPM[4317] = 12'b111111111111;
assign CPM[4318] = 12'b111111111111;
assign CPM[4319] = 12'b111111111111;
assign CPM[4320] = 12'b111111111111;
assign CPM[4321] = 12'b111111111111;
assign CPM[4322] = 12'b111111111111;
assign CPM[4323] = 12'b111111111111;
assign CPM[4324] = 12'b111111111111;
assign CPM[4325] = 12'b111111111111;
assign CPM[4326] = 12'b111111111111;
assign CPM[4327] = 12'b111111111111;
assign CPM[4328] = 12'b111111111111;
assign CPM[4329] = 12'b111111111111;
assign CPM[4330] = 12'b111111111111;
assign CPM[4331] = 12'b000000000000;
assign CPM[4332] = 12'b000000000000;
assign CPM[4333] = 12'b000000000000;
assign CPM[4334] = 12'b000000000000;
assign CPM[4335] = 12'b000000000000;
assign CPM[4336] = 12'b000000000000;
assign CPM[4337] = 12'b000000000000;
assign CPM[4338] = 12'b000000000000;
assign CPM[4339] = 12'b111111111111;
assign CPM[4340] = 12'b111111111111;
assign CPM[4341] = 12'b111111111111;
assign CPM[4342] = 12'b111111111111;
assign CPM[4343] = 12'b111111111111;
assign CPM[4344] = 12'b111111111111;
assign CPM[4345] = 12'b111111111111;
assign CPM[4346] = 12'b111111111111;
assign CPM[4347] = 12'b111111111111;
assign CPM[4348] = 12'b111111111111;
assign CPM[4349] = 12'b111111111111;
assign CPM[4350] = 12'b111111111111;
assign CPM[4351] = 12'b111111111111;
assign CPM[4352] = 12'b111111111111;
assign CPM[4353] = 12'b111111111111;
assign CPM[4354] = 12'b111111111111;
assign CPM[4355] = 12'b111111111111;
assign CPM[4356] = 12'b111111111111;
assign CPM[4357] = 12'b111111111111;
assign CPM[4358] = 12'b111111111111;
assign CPM[4359] = 12'b111111111111;
assign CPM[4360] = 12'b111111111111;
assign CPM[4361] = 12'b111111111111;
assign CPM[4362] = 12'b111111111111;
assign CPM[4363] = 12'b000000000000;
assign CPM[4364] = 12'b000000000000;
assign CPM[4365] = 12'b000000000000;
assign CPM[4366] = 12'b000000000000;
assign CPM[4367] = 12'b000000000000;
assign CPM[4368] = 12'b000000000000;
assign CPM[4369] = 12'b000000000000;
assign CPM[4370] = 12'b000000000000;
assign CPM[4371] = 12'b111111111111;
assign CPM[4372] = 12'b111111111111;
assign CPM[4373] = 12'b111111111111;
assign CPM[4374] = 12'b111111111111;
assign CPM[4375] = 12'b111111111111;
assign CPM[4376] = 12'b111111111111;
assign CPM[4377] = 12'b111111111111;
assign CPM[4378] = 12'b111111111111;
assign CPM[4379] = 12'b111111111111;
assign CPM[4380] = 12'b111111111111;
assign CPM[4381] = 12'b111111111111;
assign CPM[4382] = 12'b111111111111;
assign CPM[4383] = 12'b111111111111;
assign CPM[4384] = 12'b111111111111;
assign CPM[4385] = 12'b111111111111;
assign CPM[4386] = 12'b111111111111;
assign CPM[4387] = 12'b111111111111;
assign CPM[4388] = 12'b111111111111;
assign CPM[4389] = 12'b111111111111;
assign CPM[4390] = 12'b111111111111;
assign CPM[4391] = 12'b111111111111;
assign CPM[4392] = 12'b111111111111;
assign CPM[4393] = 12'b111111111111;
assign CPM[4394] = 12'b111111111111;
assign CPM[4395] = 12'b111111111111;
assign CPM[4396] = 12'b111111111111;
assign CPM[4397] = 12'b111111111111;
assign CPM[4398] = 12'b111111111111;
assign CPM[4399] = 12'b000000000000;
assign CPM[4400] = 12'b000000000000;
assign CPM[4401] = 12'b000000000000;
assign CPM[4402] = 12'b000000000000;
assign CPM[4403] = 12'b111111111111;
assign CPM[4404] = 12'b111111111111;
assign CPM[4405] = 12'b111111111111;
assign CPM[4406] = 12'b111111111111;
assign CPM[4407] = 12'b111111111111;
assign CPM[4408] = 12'b111111111111;
assign CPM[4409] = 12'b111111111111;
assign CPM[4410] = 12'b111111111111;
assign CPM[4411] = 12'b111111111111;
assign CPM[4412] = 12'b111111111111;
assign CPM[4413] = 12'b111111111111;
assign CPM[4414] = 12'b111111111111;
assign CPM[4415] = 12'b111111111111;
assign CPM[4416] = 12'b111111111111;
assign CPM[4417] = 12'b111111111111;
assign CPM[4418] = 12'b111111111111;
assign CPM[4419] = 12'b111111111111;
assign CPM[4420] = 12'b111111111111;
assign CPM[4421] = 12'b111111111111;
assign CPM[4422] = 12'b111111111111;
assign CPM[4423] = 12'b111111111111;
assign CPM[4424] = 12'b111111111111;
assign CPM[4425] = 12'b111111111111;
assign CPM[4426] = 12'b111111111111;
assign CPM[4427] = 12'b111111111111;
assign CPM[4428] = 12'b111111111111;
assign CPM[4429] = 12'b111111111111;
assign CPM[4430] = 12'b111111111111;
assign CPM[4431] = 12'b000000000000;
assign CPM[4432] = 12'b000000000000;
assign CPM[4433] = 12'b000000000000;
assign CPM[4434] = 12'b000000000000;
assign CPM[4435] = 12'b111111111111;
assign CPM[4436] = 12'b111111111111;
assign CPM[4437] = 12'b111111111111;
assign CPM[4438] = 12'b111111111111;
assign CPM[4439] = 12'b111111111111;
assign CPM[4440] = 12'b111111111111;
assign CPM[4441] = 12'b111111111111;
assign CPM[4442] = 12'b111111111111;
assign CPM[4443] = 12'b111111111111;
assign CPM[4444] = 12'b111111111111;
assign CPM[4445] = 12'b111111111111;
assign CPM[4446] = 12'b111111111111;
assign CPM[4447] = 12'b111111111111;
assign CPM[4448] = 12'b111111111111;
assign CPM[4449] = 12'b111111111111;
assign CPM[4450] = 12'b111111111111;
assign CPM[4451] = 12'b111111111111;
assign CPM[4452] = 12'b111111111111;
assign CPM[4453] = 12'b111111111111;
assign CPM[4454] = 12'b111111111111;
assign CPM[4455] = 12'b111111111111;
assign CPM[4456] = 12'b111111111111;
assign CPM[4457] = 12'b111111111111;
assign CPM[4458] = 12'b111111111111;
assign CPM[4459] = 12'b111111111111;
assign CPM[4460] = 12'b111111111111;
assign CPM[4461] = 12'b111111111111;
assign CPM[4462] = 12'b111111111111;
assign CPM[4463] = 12'b000000000000;
assign CPM[4464] = 12'b000000000000;
assign CPM[4465] = 12'b000000000000;
assign CPM[4466] = 12'b000000000000;
assign CPM[4467] = 12'b111111111111;
assign CPM[4468] = 12'b111111111111;
assign CPM[4469] = 12'b111111111111;
assign CPM[4470] = 12'b111111111111;
assign CPM[4471] = 12'b111111111111;
assign CPM[4472] = 12'b111111111111;
assign CPM[4473] = 12'b111111111111;
assign CPM[4474] = 12'b111111111111;
assign CPM[4475] = 12'b111111111111;
assign CPM[4476] = 12'b111111111111;
assign CPM[4477] = 12'b111111111111;
assign CPM[4478] = 12'b111111111111;
assign CPM[4479] = 12'b111111111111;
assign CPM[4480] = 12'b111111111111;
assign CPM[4481] = 12'b111111111111;
assign CPM[4482] = 12'b111111111111;
assign CPM[4483] = 12'b111111111111;
assign CPM[4484] = 12'b111111111111;
assign CPM[4485] = 12'b111111111111;
assign CPM[4486] = 12'b111111111111;
assign CPM[4487] = 12'b111111111111;
assign CPM[4488] = 12'b111111111111;
assign CPM[4489] = 12'b111111111111;
assign CPM[4490] = 12'b111111111111;
assign CPM[4491] = 12'b111111111111;
assign CPM[4492] = 12'b111111111111;
assign CPM[4493] = 12'b111111111111;
assign CPM[4494] = 12'b111111111111;
assign CPM[4495] = 12'b000000000000;
assign CPM[4496] = 12'b000000000000;
assign CPM[4497] = 12'b000000000000;
assign CPM[4498] = 12'b000000000000;
assign CPM[4499] = 12'b111111111111;
assign CPM[4500] = 12'b111111111111;
assign CPM[4501] = 12'b111111111111;
assign CPM[4502] = 12'b111111111111;
assign CPM[4503] = 12'b111111111111;
assign CPM[4504] = 12'b111111111111;
assign CPM[4505] = 12'b111111111111;
assign CPM[4506] = 12'b111111111111;
assign CPM[4507] = 12'b111111111111;
assign CPM[4508] = 12'b111111111111;
assign CPM[4509] = 12'b111111111111;
assign CPM[4510] = 12'b111111111111;
assign CPM[4511] = 12'b111111111111;
assign CPM[4512] = 12'b111111111111;
assign CPM[4513] = 12'b111111111111;
assign CPM[4514] = 12'b111111111111;
assign CPM[4515] = 12'b111111111111;
assign CPM[4516] = 12'b111111111111;
assign CPM[4517] = 12'b111111111111;
assign CPM[4518] = 12'b111111111111;
assign CPM[4519] = 12'b111111111111;
assign CPM[4520] = 12'b111111111111;
assign CPM[4521] = 12'b111111111111;
assign CPM[4522] = 12'b111111111111;
assign CPM[4523] = 12'b111111111111;
assign CPM[4524] = 12'b111111111111;
assign CPM[4525] = 12'b111111111111;
assign CPM[4526] = 12'b111111111111;
assign CPM[4527] = 12'b000000000000;
assign CPM[4528] = 12'b000000000000;
assign CPM[4529] = 12'b000000000000;
assign CPM[4530] = 12'b000000000000;
assign CPM[4531] = 12'b111111111111;
assign CPM[4532] = 12'b111111111111;
assign CPM[4533] = 12'b111111111111;
assign CPM[4534] = 12'b111111111111;
assign CPM[4535] = 12'b111111111111;
assign CPM[4536] = 12'b111111111111;
assign CPM[4537] = 12'b111111111111;
assign CPM[4538] = 12'b111111111111;
assign CPM[4539] = 12'b111111111111;
assign CPM[4540] = 12'b111111111111;
assign CPM[4541] = 12'b111111111111;
assign CPM[4542] = 12'b111111111111;
assign CPM[4543] = 12'b111111111111;
assign CPM[4544] = 12'b111111111111;
assign CPM[4545] = 12'b111111111111;
assign CPM[4546] = 12'b111111111111;
assign CPM[4547] = 12'b111111111111;
assign CPM[4548] = 12'b111111111111;
assign CPM[4549] = 12'b111111111111;
assign CPM[4550] = 12'b111111111111;
assign CPM[4551] = 12'b111111111111;
assign CPM[4552] = 12'b111111111111;
assign CPM[4553] = 12'b111111111111;
assign CPM[4554] = 12'b111111111111;
assign CPM[4555] = 12'b111111111111;
assign CPM[4556] = 12'b111111111111;
assign CPM[4557] = 12'b111111111111;
assign CPM[4558] = 12'b111111111111;
assign CPM[4559] = 12'b000000000000;
assign CPM[4560] = 12'b000000000000;
assign CPM[4561] = 12'b000000000000;
assign CPM[4562] = 12'b000000000000;
assign CPM[4563] = 12'b111111111111;
assign CPM[4564] = 12'b111111111111;
assign CPM[4565] = 12'b111111111111;
assign CPM[4566] = 12'b111111111111;
assign CPM[4567] = 12'b111111111111;
assign CPM[4568] = 12'b111111111111;
assign CPM[4569] = 12'b111111111111;
assign CPM[4570] = 12'b111111111111;
assign CPM[4571] = 12'b111111111111;
assign CPM[4572] = 12'b111111111111;
assign CPM[4573] = 12'b111111111111;
assign CPM[4574] = 12'b111111111111;
assign CPM[4575] = 12'b111111111111;
assign CPM[4576] = 12'b111111111111;
assign CPM[4577] = 12'b111111111111;
assign CPM[4578] = 12'b111111111111;
assign CPM[4579] = 12'b111111111111;
assign CPM[4580] = 12'b111111111111;
assign CPM[4581] = 12'b111111111111;
assign CPM[4582] = 12'b111111111111;
assign CPM[4583] = 12'b111111111111;
assign CPM[4584] = 12'b111111111111;
assign CPM[4585] = 12'b111111111111;
assign CPM[4586] = 12'b111111111111;
assign CPM[4587] = 12'b111111111111;
assign CPM[4588] = 12'b111111111111;
assign CPM[4589] = 12'b111111111111;
assign CPM[4590] = 12'b111111111111;
assign CPM[4591] = 12'b000000000000;
assign CPM[4592] = 12'b000000000000;
assign CPM[4593] = 12'b000000000000;
assign CPM[4594] = 12'b000000000000;
assign CPM[4595] = 12'b111111111111;
assign CPM[4596] = 12'b111111111111;
assign CPM[4597] = 12'b111111111111;
assign CPM[4598] = 12'b111111111111;
assign CPM[4599] = 12'b111111111111;
assign CPM[4600] = 12'b111111111111;
assign CPM[4601] = 12'b111111111111;
assign CPM[4602] = 12'b111111111111;
assign CPM[4603] = 12'b111111111111;
assign CPM[4604] = 12'b111111111111;
assign CPM[4605] = 12'b111111111111;
assign CPM[4606] = 12'b111111111111;
assign CPM[4607] = 12'b111111111111;
assign CPM[4608] = 12'b111111111111;
assign CPM[4609] = 12'b111111111111;
assign CPM[4610] = 12'b111111111111;
assign CPM[4611] = 12'b111111111111;
assign CPM[4612] = 12'b111111111111;
assign CPM[4613] = 12'b111111111111;
assign CPM[4614] = 12'b111111111111;
assign CPM[4615] = 12'b111111111111;
assign CPM[4616] = 12'b111111111111;
assign CPM[4617] = 12'b111111111111;
assign CPM[4618] = 12'b111111111111;
assign CPM[4619] = 12'b111111111111;
assign CPM[4620] = 12'b111111111111;
assign CPM[4621] = 12'b111111111111;
assign CPM[4622] = 12'b111111111111;
assign CPM[4623] = 12'b000000000000;
assign CPM[4624] = 12'b000000000000;
assign CPM[4625] = 12'b000000000000;
assign CPM[4626] = 12'b000000000000;
assign CPM[4627] = 12'b111111111111;
assign CPM[4628] = 12'b111111111111;
assign CPM[4629] = 12'b111111111111;
assign CPM[4630] = 12'b111111111111;
assign CPM[4631] = 12'b111111111111;
assign CPM[4632] = 12'b111111111111;
assign CPM[4633] = 12'b111111111111;
assign CPM[4634] = 12'b111111111111;
assign CPM[4635] = 12'b111111111111;
assign CPM[4636] = 12'b111111111111;
assign CPM[4637] = 12'b111111111111;
assign CPM[4638] = 12'b111111111111;
assign CPM[4639] = 12'b111111111111;
assign CPM[4640] = 12'b111111111111;
assign CPM[4641] = 12'b111111111111;
assign CPM[4642] = 12'b111111111111;
assign CPM[4643] = 12'b111111111111;
assign CPM[4644] = 12'b111111111111;
assign CPM[4645] = 12'b111111111111;
assign CPM[4646] = 12'b111111111111;
assign CPM[4647] = 12'b111111111111;
assign CPM[4648] = 12'b111111111111;
assign CPM[4649] = 12'b111111111111;
assign CPM[4650] = 12'b111111111111;
assign CPM[4651] = 12'b111111111111;
assign CPM[4652] = 12'b111111111111;
assign CPM[4653] = 12'b111111111111;
assign CPM[4654] = 12'b111111111111;
assign CPM[4655] = 12'b000000000000;
assign CPM[4656] = 12'b000000000000;
assign CPM[4657] = 12'b000000000000;
assign CPM[4658] = 12'b000000000000;
assign CPM[4659] = 12'b111111111111;
assign CPM[4660] = 12'b111111111111;
assign CPM[4661] = 12'b111111111111;
assign CPM[4662] = 12'b111111111111;
assign CPM[4663] = 12'b111111111111;
assign CPM[4664] = 12'b111111111111;
assign CPM[4665] = 12'b111111111111;
assign CPM[4666] = 12'b111111111111;
assign CPM[4667] = 12'b111111111111;
assign CPM[4668] = 12'b111111111111;
assign CPM[4669] = 12'b111111111111;
assign CPM[4670] = 12'b111111111111;
assign CPM[4671] = 12'b111111111111;
assign CPM[4672] = 12'b111111111111;
assign CPM[4673] = 12'b111111111111;
assign CPM[4674] = 12'b111111111111;
assign CPM[4675] = 12'b111111111111;
assign CPM[4676] = 12'b111111111111;
assign CPM[4677] = 12'b111111111111;
assign CPM[4678] = 12'b111111111111;
assign CPM[4679] = 12'b111111111111;
assign CPM[4680] = 12'b111111111111;
assign CPM[4681] = 12'b111111111111;
assign CPM[4682] = 12'b111111111111;
assign CPM[4683] = 12'b111111111111;
assign CPM[4684] = 12'b111111111111;
assign CPM[4685] = 12'b111111111111;
assign CPM[4686] = 12'b111111111111;
assign CPM[4687] = 12'b000000000000;
assign CPM[4688] = 12'b000000000000;
assign CPM[4689] = 12'b000000000000;
assign CPM[4690] = 12'b000000000000;
assign CPM[4691] = 12'b111111111111;
assign CPM[4692] = 12'b111111111111;
assign CPM[4693] = 12'b111111111111;
assign CPM[4694] = 12'b111111111111;
assign CPM[4695] = 12'b111111111111;
assign CPM[4696] = 12'b111111111111;
assign CPM[4697] = 12'b111111111111;
assign CPM[4698] = 12'b111111111111;
assign CPM[4699] = 12'b111111111111;
assign CPM[4700] = 12'b111111111111;
assign CPM[4701] = 12'b111111111111;
assign CPM[4702] = 12'b111111111111;
assign CPM[4703] = 12'b111111111111;
assign CPM[4704] = 12'b111111111111;
assign CPM[4705] = 12'b111111111111;
assign CPM[4706] = 12'b111111111111;
assign CPM[4707] = 12'b111111111111;
assign CPM[4708] = 12'b111111111111;
assign CPM[4709] = 12'b111111111111;
assign CPM[4710] = 12'b111111111111;
assign CPM[4711] = 12'b111111111111;
assign CPM[4712] = 12'b111111111111;
assign CPM[4713] = 12'b111111111111;
assign CPM[4714] = 12'b111111111111;
assign CPM[4715] = 12'b111111111111;
assign CPM[4716] = 12'b111111111111;
assign CPM[4717] = 12'b111111111111;
assign CPM[4718] = 12'b111111111111;
assign CPM[4719] = 12'b000000000000;
assign CPM[4720] = 12'b000000000000;
assign CPM[4721] = 12'b000000000000;
assign CPM[4722] = 12'b000000000000;
assign CPM[4723] = 12'b111111111111;
assign CPM[4724] = 12'b111111111111;
assign CPM[4725] = 12'b111111111111;
assign CPM[4726] = 12'b111111111111;
assign CPM[4727] = 12'b111111111111;
assign CPM[4728] = 12'b111111111111;
assign CPM[4729] = 12'b111111111111;
assign CPM[4730] = 12'b111111111111;
assign CPM[4731] = 12'b111111111111;
assign CPM[4732] = 12'b111111111111;
assign CPM[4733] = 12'b111111111111;
assign CPM[4734] = 12'b111111111111;
assign CPM[4735] = 12'b111111111111;
assign CPM[4736] = 12'b111111111111;
assign CPM[4737] = 12'b111111111111;
assign CPM[4738] = 12'b111111111111;
assign CPM[4739] = 12'b111111111111;
assign CPM[4740] = 12'b111111111111;
assign CPM[4741] = 12'b111111111111;
assign CPM[4742] = 12'b111111111111;
assign CPM[4743] = 12'b111111111111;
assign CPM[4744] = 12'b111111111111;
assign CPM[4745] = 12'b111111111111;
assign CPM[4746] = 12'b111111111111;
assign CPM[4747] = 12'b111111111111;
assign CPM[4748] = 12'b111111111111;
assign CPM[4749] = 12'b111111111111;
assign CPM[4750] = 12'b111111111111;
assign CPM[4751] = 12'b000000000000;
assign CPM[4752] = 12'b000000000000;
assign CPM[4753] = 12'b000000000000;
assign CPM[4754] = 12'b000000000000;
assign CPM[4755] = 12'b111111111111;
assign CPM[4756] = 12'b111111111111;
assign CPM[4757] = 12'b111111111111;
assign CPM[4758] = 12'b111111111111;
assign CPM[4759] = 12'b111111111111;
assign CPM[4760] = 12'b111111111111;
assign CPM[4761] = 12'b111111111111;
assign CPM[4762] = 12'b111111111111;
assign CPM[4763] = 12'b111111111111;
assign CPM[4764] = 12'b111111111111;
assign CPM[4765] = 12'b111111111111;
assign CPM[4766] = 12'b111111111111;
assign CPM[4767] = 12'b111111111111;
assign CPM[4768] = 12'b111111111111;
assign CPM[4769] = 12'b111111111111;
assign CPM[4770] = 12'b111111111111;
assign CPM[4771] = 12'b111111111111;
assign CPM[4772] = 12'b111111111111;
assign CPM[4773] = 12'b111111111111;
assign CPM[4774] = 12'b111111111111;
assign CPM[4775] = 12'b111111111111;
assign CPM[4776] = 12'b111111111111;
assign CPM[4777] = 12'b111111111111;
assign CPM[4778] = 12'b111111111111;
assign CPM[4779] = 12'b111111111111;
assign CPM[4780] = 12'b111111111111;
assign CPM[4781] = 12'b111111111111;
assign CPM[4782] = 12'b111111111111;
assign CPM[4783] = 12'b000000000000;
assign CPM[4784] = 12'b000000000000;
assign CPM[4785] = 12'b000000000000;
assign CPM[4786] = 12'b000000000000;
assign CPM[4787] = 12'b111111111111;
assign CPM[4788] = 12'b111111111111;
assign CPM[4789] = 12'b111111111111;
assign CPM[4790] = 12'b111111111111;
assign CPM[4791] = 12'b111111111111;
assign CPM[4792] = 12'b111111111111;
assign CPM[4793] = 12'b111111111111;
assign CPM[4794] = 12'b111111111111;
assign CPM[4795] = 12'b111111111111;
assign CPM[4796] = 12'b111111111111;
assign CPM[4797] = 12'b111111111111;
assign CPM[4798] = 12'b111111111111;
assign CPM[4799] = 12'b111111111111;
assign CPM[4800] = 12'b111111111111;
assign CPM[4801] = 12'b111111111111;
assign CPM[4802] = 12'b111111111111;
assign CPM[4803] = 12'b111111111111;
assign CPM[4804] = 12'b111111111111;
assign CPM[4805] = 12'b111111111111;
assign CPM[4806] = 12'b111111111111;
assign CPM[4807] = 12'b111111111111;
assign CPM[4808] = 12'b111111111111;
assign CPM[4809] = 12'b111111111111;
assign CPM[4810] = 12'b111111111111;
assign CPM[4811] = 12'b111111111111;
assign CPM[4812] = 12'b111111111111;
assign CPM[4813] = 12'b111111111111;
assign CPM[4814] = 12'b111111111111;
assign CPM[4815] = 12'b000000000000;
assign CPM[4816] = 12'b000000000000;
assign CPM[4817] = 12'b000000000000;
assign CPM[4818] = 12'b000000000000;
assign CPM[4819] = 12'b111111111111;
assign CPM[4820] = 12'b111111111111;
assign CPM[4821] = 12'b111111111111;
assign CPM[4822] = 12'b111111111111;
assign CPM[4823] = 12'b111111111111;
assign CPM[4824] = 12'b111111111111;
assign CPM[4825] = 12'b111111111111;
assign CPM[4826] = 12'b111111111111;
assign CPM[4827] = 12'b111111111111;
assign CPM[4828] = 12'b111111111111;
assign CPM[4829] = 12'b111111111111;
assign CPM[4830] = 12'b111111111111;
assign CPM[4831] = 12'b111111111111;
assign CPM[4832] = 12'b111111111111;
assign CPM[4833] = 12'b111111111111;
assign CPM[4834] = 12'b111111111111;
assign CPM[4835] = 12'b111111111111;
assign CPM[4836] = 12'b111111111111;
assign CPM[4837] = 12'b111111111111;
assign CPM[4838] = 12'b111111111111;
assign CPM[4839] = 12'b111111111111;
assign CPM[4840] = 12'b111111111111;
assign CPM[4841] = 12'b111111111111;
assign CPM[4842] = 12'b111111111111;
assign CPM[4843] = 12'b111111111111;
assign CPM[4844] = 12'b111111111111;
assign CPM[4845] = 12'b111111111111;
assign CPM[4846] = 12'b111111111111;
assign CPM[4847] = 12'b000000000000;
assign CPM[4848] = 12'b000000000000;
assign CPM[4849] = 12'b000000000000;
assign CPM[4850] = 12'b000000000000;
assign CPM[4851] = 12'b111111111111;
assign CPM[4852] = 12'b111111111111;
assign CPM[4853] = 12'b111111111111;
assign CPM[4854] = 12'b111111111111;
assign CPM[4855] = 12'b111111111111;
assign CPM[4856] = 12'b111111111111;
assign CPM[4857] = 12'b111111111111;
assign CPM[4858] = 12'b111111111111;
assign CPM[4859] = 12'b111111111111;
assign CPM[4860] = 12'b111111111111;
assign CPM[4861] = 12'b111111111111;
assign CPM[4862] = 12'b111111111111;
assign CPM[4863] = 12'b111111111111;
assign CPM[4864] = 12'b111111111111;
assign CPM[4865] = 12'b111111111111;
assign CPM[4866] = 12'b111111111111;
assign CPM[4867] = 12'b111111111111;
assign CPM[4868] = 12'b111111111111;
assign CPM[4869] = 12'b111111111111;
assign CPM[4870] = 12'b111111111111;
assign CPM[4871] = 12'b111111111111;
assign CPM[4872] = 12'b111111111111;
assign CPM[4873] = 12'b111111111111;
assign CPM[4874] = 12'b111111111111;
assign CPM[4875] = 12'b111111111111;
assign CPM[4876] = 12'b111111111111;
assign CPM[4877] = 12'b111111111111;
assign CPM[4878] = 12'b111111111111;
assign CPM[4879] = 12'b000000000000;
assign CPM[4880] = 12'b000000000000;
assign CPM[4881] = 12'b000000000000;
assign CPM[4882] = 12'b000000000000;
assign CPM[4883] = 12'b111111111111;
assign CPM[4884] = 12'b111111111111;
assign CPM[4885] = 12'b111111111111;
assign CPM[4886] = 12'b111111111111;
assign CPM[4887] = 12'b111111111111;
assign CPM[4888] = 12'b111111111111;
assign CPM[4889] = 12'b111111111111;
assign CPM[4890] = 12'b111111111111;
assign CPM[4891] = 12'b111111111111;
assign CPM[4892] = 12'b111111111111;
assign CPM[4893] = 12'b111111111111;
assign CPM[4894] = 12'b111111111111;
assign CPM[4895] = 12'b111111111111;
assign CPM[4896] = 12'b111111111111;
assign CPM[4897] = 12'b111111111111;
assign CPM[4898] = 12'b111111111111;
assign CPM[4899] = 12'b111111111111;
assign CPM[4900] = 12'b111111111111;
assign CPM[4901] = 12'b111111111111;
assign CPM[4902] = 12'b111111111111;
assign CPM[4903] = 12'b111111111111;
assign CPM[4904] = 12'b111111111111;
assign CPM[4905] = 12'b111111111111;
assign CPM[4906] = 12'b111111111111;
assign CPM[4907] = 12'b111111111111;
assign CPM[4908] = 12'b111111111111;
assign CPM[4909] = 12'b111111111111;
assign CPM[4910] = 12'b111111111111;
assign CPM[4911] = 12'b000000000000;
assign CPM[4912] = 12'b000000000000;
assign CPM[4913] = 12'b000000000000;
assign CPM[4914] = 12'b000000000000;
assign CPM[4915] = 12'b111111111111;
assign CPM[4916] = 12'b111111111111;
assign CPM[4917] = 12'b111111111111;
assign CPM[4918] = 12'b111111111111;
assign CPM[4919] = 12'b111111111111;
assign CPM[4920] = 12'b111111111111;
assign CPM[4921] = 12'b111111111111;
assign CPM[4922] = 12'b111111111111;
assign CPM[4923] = 12'b111111111111;
assign CPM[4924] = 12'b111111111111;
assign CPM[4925] = 12'b111111111111;
assign CPM[4926] = 12'b111111111111;
assign CPM[4927] = 12'b111111111111;
assign CPM[4928] = 12'b111111111111;
assign CPM[4929] = 12'b111111111111;
assign CPM[4930] = 12'b111111111111;
assign CPM[4931] = 12'b111111111111;
assign CPM[4932] = 12'b111111111111;
assign CPM[4933] = 12'b111111111111;
assign CPM[4934] = 12'b111111111111;
assign CPM[4935] = 12'b111111111111;
assign CPM[4936] = 12'b111111111111;
assign CPM[4937] = 12'b000000000000;
assign CPM[4938] = 12'b000000000000;
assign CPM[4939] = 12'b000000000000;
assign CPM[4940] = 12'b000000000000;
assign CPM[4941] = 12'b000000000000;
assign CPM[4942] = 12'b000000000000;
assign CPM[4943] = 12'b000000000000;
assign CPM[4944] = 12'b000000000000;
assign CPM[4945] = 12'b000000000000;
assign CPM[4946] = 12'b000000000000;
assign CPM[4947] = 12'b000000000000;
assign CPM[4948] = 12'b000000000000;
assign CPM[4949] = 12'b000000000000;
assign CPM[4950] = 12'b000000000000;
assign CPM[4951] = 12'b000000000000;
assign CPM[4952] = 12'b000000000000;
assign CPM[4953] = 12'b111111111111;
assign CPM[4954] = 12'b111111111111;
assign CPM[4955] = 12'b111111111111;
assign CPM[4956] = 12'b111111111111;
assign CPM[4957] = 12'b111111111111;
assign CPM[4958] = 12'b111111111111;
assign CPM[4959] = 12'b111111111111;
assign CPM[4960] = 12'b111111111111;
assign CPM[4961] = 12'b111111111111;
assign CPM[4962] = 12'b111111111111;
assign CPM[4963] = 12'b111111111111;
assign CPM[4964] = 12'b111111111111;
assign CPM[4965] = 12'b111111111111;
assign CPM[4966] = 12'b111111111111;
assign CPM[4967] = 12'b111111111111;
assign CPM[4968] = 12'b111111111111;
assign CPM[4969] = 12'b000000000000;
assign CPM[4970] = 12'b000000000000;
assign CPM[4971] = 12'b000000000000;
assign CPM[4972] = 12'b000000000000;
assign CPM[4973] = 12'b000000000000;
assign CPM[4974] = 12'b000000000000;
assign CPM[4975] = 12'b000000000000;
assign CPM[4976] = 12'b000000000000;
assign CPM[4977] = 12'b000000000000;
assign CPM[4978] = 12'b000000000000;
assign CPM[4979] = 12'b000000000000;
assign CPM[4980] = 12'b000000000000;
assign CPM[4981] = 12'b000000000000;
assign CPM[4982] = 12'b000000000000;
assign CPM[4983] = 12'b000000000000;
assign CPM[4984] = 12'b000000000000;
assign CPM[4985] = 12'b111111111111;
assign CPM[4986] = 12'b111111111111;
assign CPM[4987] = 12'b111111111111;
assign CPM[4988] = 12'b111111111111;
assign CPM[4989] = 12'b111111111111;
assign CPM[4990] = 12'b111111111111;
assign CPM[4991] = 12'b111111111111;
assign CPM[4992] = 12'b111111111111;
assign CPM[4993] = 12'b111111111111;
assign CPM[4994] = 12'b111111111111;
assign CPM[4995] = 12'b111111111111;
assign CPM[4996] = 12'b111111111111;
assign CPM[4997] = 12'b111111111111;
assign CPM[4998] = 12'b111111111111;
assign CPM[4999] = 12'b111111111111;
assign CPM[5000] = 12'b111111111111;
assign CPM[5001] = 12'b000000000000;
assign CPM[5002] = 12'b000000000000;
assign CPM[5003] = 12'b000000000000;
assign CPM[5004] = 12'b000000000000;
assign CPM[5005] = 12'b000000000000;
assign CPM[5006] = 12'b000000000000;
assign CPM[5007] = 12'b000000000000;
assign CPM[5008] = 12'b000000000000;
assign CPM[5009] = 12'b000000000000;
assign CPM[5010] = 12'b000000000000;
assign CPM[5011] = 12'b000000000000;
assign CPM[5012] = 12'b000000000000;
assign CPM[5013] = 12'b000000000000;
assign CPM[5014] = 12'b000000000000;
assign CPM[5015] = 12'b000000000000;
assign CPM[5016] = 12'b000000000000;
assign CPM[5017] = 12'b111111111111;
assign CPM[5018] = 12'b111111111111;
assign CPM[5019] = 12'b111111111111;
assign CPM[5020] = 12'b111111111111;
assign CPM[5021] = 12'b111111111111;
assign CPM[5022] = 12'b111111111111;
assign CPM[5023] = 12'b111111111111;
assign CPM[5024] = 12'b111111111111;
assign CPM[5025] = 12'b111111111111;
assign CPM[5026] = 12'b111111111111;
assign CPM[5027] = 12'b111111111111;
assign CPM[5028] = 12'b111111111111;
assign CPM[5029] = 12'b111111111111;
assign CPM[5030] = 12'b111111111111;
assign CPM[5031] = 12'b111111111111;
assign CPM[5032] = 12'b111111111111;
assign CPM[5033] = 12'b000000000000;
assign CPM[5034] = 12'b000000000000;
assign CPM[5035] = 12'b000000000000;
assign CPM[5036] = 12'b000000000000;
assign CPM[5037] = 12'b000000000000;
assign CPM[5038] = 12'b000000000000;
assign CPM[5039] = 12'b000000000000;
assign CPM[5040] = 12'b000000000000;
assign CPM[5041] = 12'b000000000000;
assign CPM[5042] = 12'b000000000000;
assign CPM[5043] = 12'b000000000000;
assign CPM[5044] = 12'b000000000000;
assign CPM[5045] = 12'b000000000000;
assign CPM[5046] = 12'b000000000000;
assign CPM[5047] = 12'b000000000000;
assign CPM[5048] = 12'b000000000000;
assign CPM[5049] = 12'b111111111111;
assign CPM[5050] = 12'b111111111111;
assign CPM[5051] = 12'b111111111111;
assign CPM[5052] = 12'b111111111111;
assign CPM[5053] = 12'b111111111111;
assign CPM[5054] = 12'b111111111111;
assign CPM[5055] = 12'b111111111111;
assign CPM[5056] = 12'b111111111111;
assign CPM[5057] = 12'b111111111111;
assign CPM[5058] = 12'b111111111111;
assign CPM[5059] = 12'b111111111111;
assign CPM[5060] = 12'b111111111111;
assign CPM[5061] = 12'b111111111111;
assign CPM[5062] = 12'b111111111111;
assign CPM[5063] = 12'b111111111111;
assign CPM[5064] = 12'b111111111111;
assign CPM[5065] = 12'b111111111111;
assign CPM[5066] = 12'b111111111111;
assign CPM[5067] = 12'b111111111111;
assign CPM[5068] = 12'b111111111111;
assign CPM[5069] = 12'b111111111111;
assign CPM[5070] = 12'b111111111111;
assign CPM[5071] = 12'b111111111111;
assign CPM[5072] = 12'b111111111111;
assign CPM[5073] = 12'b111111111111;
assign CPM[5074] = 12'b111111111111;
assign CPM[5075] = 12'b111111111111;
assign CPM[5076] = 12'b111111111111;
assign CPM[5077] = 12'b111111111111;
assign CPM[5078] = 12'b111111111111;
assign CPM[5079] = 12'b111111111111;
assign CPM[5080] = 12'b111111111111;
assign CPM[5081] = 12'b111111111111;
assign CPM[5082] = 12'b111111111111;
assign CPM[5083] = 12'b111111111111;
assign CPM[5084] = 12'b111111111111;
assign CPM[5085] = 12'b111111111111;
assign CPM[5086] = 12'b111111111111;
assign CPM[5087] = 12'b111111111111;
assign CPM[5088] = 12'b111111111111;
assign CPM[5089] = 12'b111111111111;
assign CPM[5090] = 12'b111111111111;
assign CPM[5091] = 12'b111111111111;
assign CPM[5092] = 12'b111111111111;
assign CPM[5093] = 12'b111111111111;
assign CPM[5094] = 12'b111111111111;
assign CPM[5095] = 12'b111111111111;
assign CPM[5096] = 12'b111111111111;
assign CPM[5097] = 12'b111111111111;
assign CPM[5098] = 12'b111111111111;
assign CPM[5099] = 12'b111111111111;
assign CPM[5100] = 12'b111111111111;
assign CPM[5101] = 12'b111111111111;
assign CPM[5102] = 12'b111111111111;
assign CPM[5103] = 12'b111111111111;
assign CPM[5104] = 12'b111111111111;
assign CPM[5105] = 12'b111111111111;
assign CPM[5106] = 12'b111111111111;
assign CPM[5107] = 12'b111111111111;
assign CPM[5108] = 12'b111111111111;
assign CPM[5109] = 12'b111111111111;
assign CPM[5110] = 12'b111111111111;
assign CPM[5111] = 12'b111111111111;
assign CPM[5112] = 12'b111111111111;
assign CPM[5113] = 12'b111111111111;
assign CPM[5114] = 12'b111111111111;
assign CPM[5115] = 12'b111111111111;
assign CPM[5116] = 12'b111111111111;
assign CPM[5117] = 12'b111111111111;
assign CPM[5118] = 12'b111111111111;
assign CPM[5119] = 12'b111111111111;
assign CPM[5120] = 12'b111111111111;
assign CPM[5121] = 12'b111111111111;
assign CPM[5122] = 12'b111111111111;
assign CPM[5123] = 12'b111111111111;
assign CPM[5124] = 12'b111111111111;
assign CPM[5125] = 12'b111111111111;
assign CPM[5126] = 12'b111111111111;
assign CPM[5127] = 12'b111111111111;
assign CPM[5128] = 12'b111111111111;
assign CPM[5129] = 12'b111111111111;
assign CPM[5130] = 12'b111111111111;
assign CPM[5131] = 12'b111111111111;
assign CPM[5132] = 12'b111111111111;
assign CPM[5133] = 12'b111111111111;
assign CPM[5134] = 12'b111111111111;
assign CPM[5135] = 12'b111111111111;
assign CPM[5136] = 12'b111111111111;
assign CPM[5137] = 12'b111111111111;
assign CPM[5138] = 12'b111111111111;
assign CPM[5139] = 12'b111111111111;
assign CPM[5140] = 12'b111111111111;
assign CPM[5141] = 12'b111111111111;
assign CPM[5142] = 12'b111111111111;
assign CPM[5143] = 12'b111111111111;
assign CPM[5144] = 12'b111111111111;
assign CPM[5145] = 12'b111111111111;
assign CPM[5146] = 12'b111111111111;
assign CPM[5147] = 12'b111111111111;
assign CPM[5148] = 12'b111111111111;
assign CPM[5149] = 12'b111111111111;
assign CPM[5150] = 12'b111111111111;
assign CPM[5151] = 12'b111111111111;
assign CPM[5152] = 12'b111111111111;
assign CPM[5153] = 12'b111111111111;
assign CPM[5154] = 12'b111111111111;
assign CPM[5155] = 12'b111111111111;
assign CPM[5156] = 12'b111111111111;
assign CPM[5157] = 12'b111111111111;
assign CPM[5158] = 12'b111111111111;
assign CPM[5159] = 12'b111111111111;
assign CPM[5160] = 12'b111111111111;
assign CPM[5161] = 12'b111111111111;
assign CPM[5162] = 12'b111111111111;
assign CPM[5163] = 12'b111111111111;
assign CPM[5164] = 12'b111111111111;
assign CPM[5165] = 12'b111111111111;
assign CPM[5166] = 12'b111111111111;
assign CPM[5167] = 12'b111111111111;
assign CPM[5168] = 12'b111111111111;
assign CPM[5169] = 12'b111111111111;
assign CPM[5170] = 12'b111111111111;
assign CPM[5171] = 12'b111111111111;
assign CPM[5172] = 12'b111111111111;
assign CPM[5173] = 12'b111111111111;
assign CPM[5174] = 12'b111111111111;
assign CPM[5175] = 12'b111111111111;
assign CPM[5176] = 12'b111111111111;
assign CPM[5177] = 12'b111111111111;
assign CPM[5178] = 12'b111111111111;
assign CPM[5179] = 12'b111111111111;
assign CPM[5180] = 12'b111111111111;
assign CPM[5181] = 12'b111111111111;
assign CPM[5182] = 12'b111111111111;
assign CPM[5183] = 12'b111111111111;
assign CPM[5184] = 12'b111111111111;
assign CPM[5185] = 12'b111111111111;
assign CPM[5186] = 12'b111111111111;
assign CPM[5187] = 12'b111111111111;
assign CPM[5188] = 12'b111111111111;
assign CPM[5189] = 12'b111111111111;
assign CPM[5190] = 12'b111111111111;
assign CPM[5191] = 12'b111111111111;
assign CPM[5192] = 12'b111111111111;
assign CPM[5193] = 12'b111111111111;
assign CPM[5194] = 12'b111111111111;
assign CPM[5195] = 12'b111111111111;
assign CPM[5196] = 12'b111111111111;
assign CPM[5197] = 12'b111111111111;
assign CPM[5198] = 12'b111111111111;
assign CPM[5199] = 12'b111111111111;
assign CPM[5200] = 12'b111111111111;
assign CPM[5201] = 12'b111111111111;
assign CPM[5202] = 12'b111111111111;
assign CPM[5203] = 12'b111111111111;
assign CPM[5204] = 12'b111111111111;
assign CPM[5205] = 12'b111111111111;
assign CPM[5206] = 12'b111111111111;
assign CPM[5207] = 12'b111111111111;
assign CPM[5208] = 12'b111111111111;
assign CPM[5209] = 12'b111111111111;
assign CPM[5210] = 12'b111111111111;
assign CPM[5211] = 12'b111111111111;
assign CPM[5212] = 12'b111111111111;
assign CPM[5213] = 12'b111111111111;
assign CPM[5214] = 12'b111111111111;
assign CPM[5215] = 12'b111111111111;
assign CPM[5216] = 12'b111111111111;
assign CPM[5217] = 12'b111111111111;
assign CPM[5218] = 12'b111111111111;
assign CPM[5219] = 12'b111111111111;
assign CPM[5220] = 12'b111111111111;
assign CPM[5221] = 12'b111111111111;
assign CPM[5222] = 12'b111111111111;
assign CPM[5223] = 12'b111111111111;
assign CPM[5224] = 12'b111111111111;
assign CPM[5225] = 12'b111111111111;
assign CPM[5226] = 12'b111111111111;
assign CPM[5227] = 12'b111111111111;
assign CPM[5228] = 12'b111111111111;
assign CPM[5229] = 12'b111111111111;
assign CPM[5230] = 12'b111111111111;
assign CPM[5231] = 12'b111111111111;
assign CPM[5232] = 12'b111111111111;
assign CPM[5233] = 12'b111111111111;
assign CPM[5234] = 12'b111111111111;
assign CPM[5235] = 12'b111111111111;
assign CPM[5236] = 12'b111111111111;
assign CPM[5237] = 12'b111111111111;
assign CPM[5238] = 12'b111111111111;
assign CPM[5239] = 12'b111111111111;
assign CPM[5240] = 12'b111111111111;
assign CPM[5241] = 12'b111111111111;
assign CPM[5242] = 12'b111111111111;
assign CPM[5243] = 12'b111111111111;
assign CPM[5244] = 12'b111111111111;
assign CPM[5245] = 12'b111111111111;
assign CPM[5246] = 12'b111111111111;
assign CPM[5247] = 12'b111111111111;
assign CPM[5248] = 12'b111111111111;
assign CPM[5249] = 12'b111111111111;
assign CPM[5250] = 12'b111111111111;
assign CPM[5251] = 12'b111111111111;
assign CPM[5252] = 12'b111111111111;
assign CPM[5253] = 12'b111111111111;
assign CPM[5254] = 12'b111111111111;
assign CPM[5255] = 12'b111111111111;
assign CPM[5256] = 12'b111111111111;
assign CPM[5257] = 12'b111111111111;
assign CPM[5258] = 12'b111111111111;
assign CPM[5259] = 12'b000000000000;
assign CPM[5260] = 12'b000000000000;
assign CPM[5261] = 12'b000000000000;
assign CPM[5262] = 12'b000000000000;
assign CPM[5263] = 12'b000000000000;
assign CPM[5264] = 12'b000000000000;
assign CPM[5265] = 12'b000000000000;
assign CPM[5266] = 12'b000000000000;
assign CPM[5267] = 12'b000000000000;
assign CPM[5268] = 12'b000000000000;
assign CPM[5269] = 12'b111111111111;
assign CPM[5270] = 12'b111111111111;
assign CPM[5271] = 12'b111111111111;
assign CPM[5272] = 12'b111111111111;
assign CPM[5273] = 12'b111111111111;
assign CPM[5274] = 12'b111111111111;
assign CPM[5275] = 12'b111111111111;
assign CPM[5276] = 12'b111111111111;
assign CPM[5277] = 12'b111111111111;
assign CPM[5278] = 12'b111111111111;
assign CPM[5279] = 12'b111111111111;
assign CPM[5280] = 12'b111111111111;
assign CPM[5281] = 12'b111111111111;
assign CPM[5282] = 12'b111111111111;
assign CPM[5283] = 12'b111111111111;
assign CPM[5284] = 12'b111111111111;
assign CPM[5285] = 12'b111111111111;
assign CPM[5286] = 12'b111111111111;
assign CPM[5287] = 12'b111111111111;
assign CPM[5288] = 12'b111111111111;
assign CPM[5289] = 12'b111111111111;
assign CPM[5290] = 12'b111111111111;
assign CPM[5291] = 12'b000000000000;
assign CPM[5292] = 12'b000000000000;
assign CPM[5293] = 12'b000000000000;
assign CPM[5294] = 12'b000000000000;
assign CPM[5295] = 12'b000000000000;
assign CPM[5296] = 12'b000000000000;
assign CPM[5297] = 12'b000000000000;
assign CPM[5298] = 12'b000000000000;
assign CPM[5299] = 12'b000000000000;
assign CPM[5300] = 12'b000000000000;
assign CPM[5301] = 12'b111111111111;
assign CPM[5302] = 12'b111111111111;
assign CPM[5303] = 12'b111111111111;
assign CPM[5304] = 12'b111111111111;
assign CPM[5305] = 12'b111111111111;
assign CPM[5306] = 12'b111111111111;
assign CPM[5307] = 12'b111111111111;
assign CPM[5308] = 12'b111111111111;
assign CPM[5309] = 12'b111111111111;
assign CPM[5310] = 12'b111111111111;
assign CPM[5311] = 12'b111111111111;
assign CPM[5312] = 12'b111111111111;
assign CPM[5313] = 12'b111111111111;
assign CPM[5314] = 12'b111111111111;
assign CPM[5315] = 12'b111111111111;
assign CPM[5316] = 12'b111111111111;
assign CPM[5317] = 12'b111111111111;
assign CPM[5318] = 12'b111111111111;
assign CPM[5319] = 12'b111111111111;
assign CPM[5320] = 12'b111111111111;
assign CPM[5321] = 12'b111111111111;
assign CPM[5322] = 12'b111111111111;
assign CPM[5323] = 12'b000000000000;
assign CPM[5324] = 12'b000000000000;
assign CPM[5325] = 12'b000000000000;
assign CPM[5326] = 12'b000000000000;
assign CPM[5327] = 12'b000000000000;
assign CPM[5328] = 12'b000000000000;
assign CPM[5329] = 12'b000000000000;
assign CPM[5330] = 12'b000000000000;
assign CPM[5331] = 12'b000000000000;
assign CPM[5332] = 12'b000000000000;
assign CPM[5333] = 12'b111111111111;
assign CPM[5334] = 12'b111111111111;
assign CPM[5335] = 12'b111111111111;
assign CPM[5336] = 12'b111111111111;
assign CPM[5337] = 12'b111111111111;
assign CPM[5338] = 12'b111111111111;
assign CPM[5339] = 12'b111111111111;
assign CPM[5340] = 12'b111111111111;
assign CPM[5341] = 12'b111111111111;
assign CPM[5342] = 12'b111111111111;
assign CPM[5343] = 12'b111111111111;
assign CPM[5344] = 12'b111111111111;
assign CPM[5345] = 12'b111111111111;
assign CPM[5346] = 12'b111111111111;
assign CPM[5347] = 12'b111111111111;
assign CPM[5348] = 12'b111111111111;
assign CPM[5349] = 12'b111111111111;
assign CPM[5350] = 12'b111111111111;
assign CPM[5351] = 12'b111111111111;
assign CPM[5352] = 12'b111111111111;
assign CPM[5353] = 12'b111111111111;
assign CPM[5354] = 12'b111111111111;
assign CPM[5355] = 12'b000000000000;
assign CPM[5356] = 12'b000000000000;
assign CPM[5357] = 12'b000000000000;
assign CPM[5358] = 12'b000000000000;
assign CPM[5359] = 12'b000000000000;
assign CPM[5360] = 12'b000000000000;
assign CPM[5361] = 12'b000000000000;
assign CPM[5362] = 12'b000000000000;
assign CPM[5363] = 12'b000000000000;
assign CPM[5364] = 12'b000000000000;
assign CPM[5365] = 12'b111111111111;
assign CPM[5366] = 12'b111111111111;
assign CPM[5367] = 12'b111111111111;
assign CPM[5368] = 12'b111111111111;
assign CPM[5369] = 12'b111111111111;
assign CPM[5370] = 12'b111111111111;
assign CPM[5371] = 12'b111111111111;
assign CPM[5372] = 12'b111111111111;
assign CPM[5373] = 12'b111111111111;
assign CPM[5374] = 12'b111111111111;
assign CPM[5375] = 12'b111111111111;
assign CPM[5376] = 12'b111111111111;
assign CPM[5377] = 12'b111111111111;
assign CPM[5378] = 12'b111111111111;
assign CPM[5379] = 12'b111111111111;
assign CPM[5380] = 12'b111111111111;
assign CPM[5381] = 12'b111111111111;
assign CPM[5382] = 12'b111111111111;
assign CPM[5383] = 12'b000000000000;
assign CPM[5384] = 12'b000000000000;
assign CPM[5385] = 12'b000000000000;
assign CPM[5386] = 12'b000000000000;
assign CPM[5387] = 12'b111111111111;
assign CPM[5388] = 12'b111111111111;
assign CPM[5389] = 12'b111111111111;
assign CPM[5390] = 12'b111111111111;
assign CPM[5391] = 12'b111111111111;
assign CPM[5392] = 12'b111111111111;
assign CPM[5393] = 12'b111111111111;
assign CPM[5394] = 12'b111111111111;
assign CPM[5395] = 12'b111111111111;
assign CPM[5396] = 12'b111111111111;
assign CPM[5397] = 12'b000000000000;
assign CPM[5398] = 12'b000000000000;
assign CPM[5399] = 12'b000000000000;
assign CPM[5400] = 12'b000000000000;
assign CPM[5401] = 12'b111111111111;
assign CPM[5402] = 12'b111111111111;
assign CPM[5403] = 12'b111111111111;
assign CPM[5404] = 12'b111111111111;
assign CPM[5405] = 12'b111111111111;
assign CPM[5406] = 12'b111111111111;
assign CPM[5407] = 12'b111111111111;
assign CPM[5408] = 12'b111111111111;
assign CPM[5409] = 12'b111111111111;
assign CPM[5410] = 12'b111111111111;
assign CPM[5411] = 12'b111111111111;
assign CPM[5412] = 12'b111111111111;
assign CPM[5413] = 12'b111111111111;
assign CPM[5414] = 12'b111111111111;
assign CPM[5415] = 12'b000000000000;
assign CPM[5416] = 12'b000000000000;
assign CPM[5417] = 12'b000000000000;
assign CPM[5418] = 12'b000000000000;
assign CPM[5419] = 12'b111111111111;
assign CPM[5420] = 12'b111111111111;
assign CPM[5421] = 12'b111111111111;
assign CPM[5422] = 12'b111111111111;
assign CPM[5423] = 12'b111111111111;
assign CPM[5424] = 12'b111111111111;
assign CPM[5425] = 12'b111111111111;
assign CPM[5426] = 12'b111111111111;
assign CPM[5427] = 12'b111111111111;
assign CPM[5428] = 12'b111111111111;
assign CPM[5429] = 12'b000000000000;
assign CPM[5430] = 12'b000000000000;
assign CPM[5431] = 12'b000000000000;
assign CPM[5432] = 12'b000000000000;
assign CPM[5433] = 12'b111111111111;
assign CPM[5434] = 12'b111111111111;
assign CPM[5435] = 12'b111111111111;
assign CPM[5436] = 12'b111111111111;
assign CPM[5437] = 12'b111111111111;
assign CPM[5438] = 12'b111111111111;
assign CPM[5439] = 12'b111111111111;
assign CPM[5440] = 12'b111111111111;
assign CPM[5441] = 12'b111111111111;
assign CPM[5442] = 12'b111111111111;
assign CPM[5443] = 12'b111111111111;
assign CPM[5444] = 12'b111111111111;
assign CPM[5445] = 12'b111111111111;
assign CPM[5446] = 12'b111111111111;
assign CPM[5447] = 12'b000000000000;
assign CPM[5448] = 12'b000000000000;
assign CPM[5449] = 12'b000000000000;
assign CPM[5450] = 12'b000000000000;
assign CPM[5451] = 12'b111111111111;
assign CPM[5452] = 12'b111111111111;
assign CPM[5453] = 12'b111111111111;
assign CPM[5454] = 12'b111111111111;
assign CPM[5455] = 12'b111111111111;
assign CPM[5456] = 12'b111111111111;
assign CPM[5457] = 12'b111111111111;
assign CPM[5458] = 12'b111111111111;
assign CPM[5459] = 12'b111111111111;
assign CPM[5460] = 12'b111111111111;
assign CPM[5461] = 12'b000000000000;
assign CPM[5462] = 12'b000000000000;
assign CPM[5463] = 12'b000000000000;
assign CPM[5464] = 12'b000000000000;
assign CPM[5465] = 12'b111111111111;
assign CPM[5466] = 12'b111111111111;
assign CPM[5467] = 12'b111111111111;
assign CPM[5468] = 12'b111111111111;
assign CPM[5469] = 12'b111111111111;
assign CPM[5470] = 12'b111111111111;
assign CPM[5471] = 12'b111111111111;
assign CPM[5472] = 12'b111111111111;
assign CPM[5473] = 12'b111111111111;
assign CPM[5474] = 12'b111111111111;
assign CPM[5475] = 12'b111111111111;
assign CPM[5476] = 12'b111111111111;
assign CPM[5477] = 12'b111111111111;
assign CPM[5478] = 12'b111111111111;
assign CPM[5479] = 12'b000000000000;
assign CPM[5480] = 12'b000000000000;
assign CPM[5481] = 12'b000000000000;
assign CPM[5482] = 12'b000000000000;
assign CPM[5483] = 12'b111111111111;
assign CPM[5484] = 12'b111111111111;
assign CPM[5485] = 12'b111111111111;
assign CPM[5486] = 12'b111111111111;
assign CPM[5487] = 12'b111111111111;
assign CPM[5488] = 12'b111111111111;
assign CPM[5489] = 12'b111111111111;
assign CPM[5490] = 12'b111111111111;
assign CPM[5491] = 12'b111111111111;
assign CPM[5492] = 12'b111111111111;
assign CPM[5493] = 12'b000000000000;
assign CPM[5494] = 12'b000000000000;
assign CPM[5495] = 12'b000000000000;
assign CPM[5496] = 12'b000000000000;
assign CPM[5497] = 12'b111111111111;
assign CPM[5498] = 12'b111111111111;
assign CPM[5499] = 12'b111111111111;
assign CPM[5500] = 12'b111111111111;
assign CPM[5501] = 12'b111111111111;
assign CPM[5502] = 12'b111111111111;
assign CPM[5503] = 12'b111111111111;
assign CPM[5504] = 12'b111111111111;
assign CPM[5505] = 12'b111111111111;
assign CPM[5506] = 12'b111111111111;
assign CPM[5507] = 12'b111111111111;
assign CPM[5508] = 12'b111111111111;
assign CPM[5509] = 12'b111111111111;
assign CPM[5510] = 12'b111111111111;
assign CPM[5511] = 12'b111111111111;
assign CPM[5512] = 12'b111111111111;
assign CPM[5513] = 12'b111111111111;
assign CPM[5514] = 12'b111111111111;
assign CPM[5515] = 12'b111111111111;
assign CPM[5516] = 12'b111111111111;
assign CPM[5517] = 12'b111111111111;
assign CPM[5518] = 12'b111111111111;
assign CPM[5519] = 12'b111111111111;
assign CPM[5520] = 12'b111111111111;
assign CPM[5521] = 12'b000000000000;
assign CPM[5522] = 12'b000000000000;
assign CPM[5523] = 12'b000000000000;
assign CPM[5524] = 12'b000000000000;
assign CPM[5525] = 12'b111111111111;
assign CPM[5526] = 12'b111111111111;
assign CPM[5527] = 12'b111111111111;
assign CPM[5528] = 12'b111111111111;
assign CPM[5529] = 12'b111111111111;
assign CPM[5530] = 12'b111111111111;
assign CPM[5531] = 12'b111111111111;
assign CPM[5532] = 12'b111111111111;
assign CPM[5533] = 12'b111111111111;
assign CPM[5534] = 12'b111111111111;
assign CPM[5535] = 12'b111111111111;
assign CPM[5536] = 12'b111111111111;
assign CPM[5537] = 12'b111111111111;
assign CPM[5538] = 12'b111111111111;
assign CPM[5539] = 12'b111111111111;
assign CPM[5540] = 12'b111111111111;
assign CPM[5541] = 12'b111111111111;
assign CPM[5542] = 12'b111111111111;
assign CPM[5543] = 12'b111111111111;
assign CPM[5544] = 12'b111111111111;
assign CPM[5545] = 12'b111111111111;
assign CPM[5546] = 12'b111111111111;
assign CPM[5547] = 12'b111111111111;
assign CPM[5548] = 12'b111111111111;
assign CPM[5549] = 12'b111111111111;
assign CPM[5550] = 12'b111111111111;
assign CPM[5551] = 12'b111111111111;
assign CPM[5552] = 12'b111111111111;
assign CPM[5553] = 12'b000000000000;
assign CPM[5554] = 12'b000000000000;
assign CPM[5555] = 12'b000000000000;
assign CPM[5556] = 12'b000000000000;
assign CPM[5557] = 12'b111111111111;
assign CPM[5558] = 12'b111111111111;
assign CPM[5559] = 12'b111111111111;
assign CPM[5560] = 12'b111111111111;
assign CPM[5561] = 12'b111111111111;
assign CPM[5562] = 12'b111111111111;
assign CPM[5563] = 12'b111111111111;
assign CPM[5564] = 12'b111111111111;
assign CPM[5565] = 12'b111111111111;
assign CPM[5566] = 12'b111111111111;
assign CPM[5567] = 12'b111111111111;
assign CPM[5568] = 12'b111111111111;
assign CPM[5569] = 12'b111111111111;
assign CPM[5570] = 12'b111111111111;
assign CPM[5571] = 12'b111111111111;
assign CPM[5572] = 12'b111111111111;
assign CPM[5573] = 12'b111111111111;
assign CPM[5574] = 12'b111111111111;
assign CPM[5575] = 12'b111111111111;
assign CPM[5576] = 12'b111111111111;
assign CPM[5577] = 12'b111111111111;
assign CPM[5578] = 12'b111111111111;
assign CPM[5579] = 12'b111111111111;
assign CPM[5580] = 12'b111111111111;
assign CPM[5581] = 12'b111111111111;
assign CPM[5582] = 12'b111111111111;
assign CPM[5583] = 12'b111111111111;
assign CPM[5584] = 12'b111111111111;
assign CPM[5585] = 12'b000000000000;
assign CPM[5586] = 12'b000000000000;
assign CPM[5587] = 12'b000000000000;
assign CPM[5588] = 12'b000000000000;
assign CPM[5589] = 12'b111111111111;
assign CPM[5590] = 12'b111111111111;
assign CPM[5591] = 12'b111111111111;
assign CPM[5592] = 12'b111111111111;
assign CPM[5593] = 12'b111111111111;
assign CPM[5594] = 12'b111111111111;
assign CPM[5595] = 12'b111111111111;
assign CPM[5596] = 12'b111111111111;
assign CPM[5597] = 12'b111111111111;
assign CPM[5598] = 12'b111111111111;
assign CPM[5599] = 12'b111111111111;
assign CPM[5600] = 12'b111111111111;
assign CPM[5601] = 12'b111111111111;
assign CPM[5602] = 12'b111111111111;
assign CPM[5603] = 12'b111111111111;
assign CPM[5604] = 12'b111111111111;
assign CPM[5605] = 12'b111111111111;
assign CPM[5606] = 12'b111111111111;
assign CPM[5607] = 12'b111111111111;
assign CPM[5608] = 12'b111111111111;
assign CPM[5609] = 12'b111111111111;
assign CPM[5610] = 12'b111111111111;
assign CPM[5611] = 12'b111111111111;
assign CPM[5612] = 12'b111111111111;
assign CPM[5613] = 12'b111111111111;
assign CPM[5614] = 12'b111111111111;
assign CPM[5615] = 12'b111111111111;
assign CPM[5616] = 12'b111111111111;
assign CPM[5617] = 12'b000000000000;
assign CPM[5618] = 12'b000000000000;
assign CPM[5619] = 12'b000000000000;
assign CPM[5620] = 12'b000000000000;
assign CPM[5621] = 12'b111111111111;
assign CPM[5622] = 12'b111111111111;
assign CPM[5623] = 12'b111111111111;
assign CPM[5624] = 12'b111111111111;
assign CPM[5625] = 12'b111111111111;
assign CPM[5626] = 12'b111111111111;
assign CPM[5627] = 12'b111111111111;
assign CPM[5628] = 12'b111111111111;
assign CPM[5629] = 12'b111111111111;
assign CPM[5630] = 12'b111111111111;
assign CPM[5631] = 12'b111111111111;
assign CPM[5632] = 12'b111111111111;
assign CPM[5633] = 12'b111111111111;
assign CPM[5634] = 12'b111111111111;
assign CPM[5635] = 12'b111111111111;
assign CPM[5636] = 12'b111111111111;
assign CPM[5637] = 12'b111111111111;
assign CPM[5638] = 12'b111111111111;
assign CPM[5639] = 12'b111111111111;
assign CPM[5640] = 12'b111111111111;
assign CPM[5641] = 12'b111111111111;
assign CPM[5642] = 12'b111111111111;
assign CPM[5643] = 12'b111111111111;
assign CPM[5644] = 12'b111111111111;
assign CPM[5645] = 12'b000000000000;
assign CPM[5646] = 12'b000000000000;
assign CPM[5647] = 12'b000000000000;
assign CPM[5648] = 12'b000000000000;
assign CPM[5649] = 12'b111111111111;
assign CPM[5650] = 12'b111111111111;
assign CPM[5651] = 12'b111111111111;
assign CPM[5652] = 12'b111111111111;
assign CPM[5653] = 12'b111111111111;
assign CPM[5654] = 12'b111111111111;
assign CPM[5655] = 12'b111111111111;
assign CPM[5656] = 12'b111111111111;
assign CPM[5657] = 12'b111111111111;
assign CPM[5658] = 12'b111111111111;
assign CPM[5659] = 12'b111111111111;
assign CPM[5660] = 12'b111111111111;
assign CPM[5661] = 12'b111111111111;
assign CPM[5662] = 12'b111111111111;
assign CPM[5663] = 12'b111111111111;
assign CPM[5664] = 12'b111111111111;
assign CPM[5665] = 12'b111111111111;
assign CPM[5666] = 12'b111111111111;
assign CPM[5667] = 12'b111111111111;
assign CPM[5668] = 12'b111111111111;
assign CPM[5669] = 12'b111111111111;
assign CPM[5670] = 12'b111111111111;
assign CPM[5671] = 12'b111111111111;
assign CPM[5672] = 12'b111111111111;
assign CPM[5673] = 12'b111111111111;
assign CPM[5674] = 12'b111111111111;
assign CPM[5675] = 12'b111111111111;
assign CPM[5676] = 12'b111111111111;
assign CPM[5677] = 12'b000000000000;
assign CPM[5678] = 12'b000000000000;
assign CPM[5679] = 12'b000000000000;
assign CPM[5680] = 12'b000000000000;
assign CPM[5681] = 12'b111111111111;
assign CPM[5682] = 12'b111111111111;
assign CPM[5683] = 12'b111111111111;
assign CPM[5684] = 12'b111111111111;
assign CPM[5685] = 12'b111111111111;
assign CPM[5686] = 12'b111111111111;
assign CPM[5687] = 12'b111111111111;
assign CPM[5688] = 12'b111111111111;
assign CPM[5689] = 12'b111111111111;
assign CPM[5690] = 12'b111111111111;
assign CPM[5691] = 12'b111111111111;
assign CPM[5692] = 12'b111111111111;
assign CPM[5693] = 12'b111111111111;
assign CPM[5694] = 12'b111111111111;
assign CPM[5695] = 12'b111111111111;
assign CPM[5696] = 12'b111111111111;
assign CPM[5697] = 12'b111111111111;
assign CPM[5698] = 12'b111111111111;
assign CPM[5699] = 12'b111111111111;
assign CPM[5700] = 12'b111111111111;
assign CPM[5701] = 12'b111111111111;
assign CPM[5702] = 12'b111111111111;
assign CPM[5703] = 12'b111111111111;
assign CPM[5704] = 12'b111111111111;
assign CPM[5705] = 12'b111111111111;
assign CPM[5706] = 12'b111111111111;
assign CPM[5707] = 12'b111111111111;
assign CPM[5708] = 12'b111111111111;
assign CPM[5709] = 12'b000000000000;
assign CPM[5710] = 12'b000000000000;
assign CPM[5711] = 12'b000000000000;
assign CPM[5712] = 12'b000000000000;
assign CPM[5713] = 12'b111111111111;
assign CPM[5714] = 12'b111111111111;
assign CPM[5715] = 12'b111111111111;
assign CPM[5716] = 12'b111111111111;
assign CPM[5717] = 12'b111111111111;
assign CPM[5718] = 12'b111111111111;
assign CPM[5719] = 12'b111111111111;
assign CPM[5720] = 12'b111111111111;
assign CPM[5721] = 12'b111111111111;
assign CPM[5722] = 12'b111111111111;
assign CPM[5723] = 12'b111111111111;
assign CPM[5724] = 12'b111111111111;
assign CPM[5725] = 12'b111111111111;
assign CPM[5726] = 12'b111111111111;
assign CPM[5727] = 12'b111111111111;
assign CPM[5728] = 12'b111111111111;
assign CPM[5729] = 12'b111111111111;
assign CPM[5730] = 12'b111111111111;
assign CPM[5731] = 12'b111111111111;
assign CPM[5732] = 12'b111111111111;
assign CPM[5733] = 12'b111111111111;
assign CPM[5734] = 12'b111111111111;
assign CPM[5735] = 12'b111111111111;
assign CPM[5736] = 12'b111111111111;
assign CPM[5737] = 12'b111111111111;
assign CPM[5738] = 12'b111111111111;
assign CPM[5739] = 12'b111111111111;
assign CPM[5740] = 12'b111111111111;
assign CPM[5741] = 12'b000000000000;
assign CPM[5742] = 12'b000000000000;
assign CPM[5743] = 12'b000000000000;
assign CPM[5744] = 12'b000000000000;
assign CPM[5745] = 12'b111111111111;
assign CPM[5746] = 12'b111111111111;
assign CPM[5747] = 12'b111111111111;
assign CPM[5748] = 12'b111111111111;
assign CPM[5749] = 12'b111111111111;
assign CPM[5750] = 12'b111111111111;
assign CPM[5751] = 12'b111111111111;
assign CPM[5752] = 12'b111111111111;
assign CPM[5753] = 12'b111111111111;
assign CPM[5754] = 12'b111111111111;
assign CPM[5755] = 12'b111111111111;
assign CPM[5756] = 12'b111111111111;
assign CPM[5757] = 12'b111111111111;
assign CPM[5758] = 12'b111111111111;
assign CPM[5759] = 12'b111111111111;
assign CPM[5760] = 12'b111111111111;
assign CPM[5761] = 12'b111111111111;
assign CPM[5762] = 12'b111111111111;
assign CPM[5763] = 12'b111111111111;
assign CPM[5764] = 12'b111111111111;
assign CPM[5765] = 12'b111111111111;
assign CPM[5766] = 12'b111111111111;
assign CPM[5767] = 12'b111111111111;
assign CPM[5768] = 12'b111111111111;
assign CPM[5769] = 12'b000000000000;
assign CPM[5770] = 12'b000000000000;
assign CPM[5771] = 12'b000000000000;
assign CPM[5772] = 12'b000000000000;
assign CPM[5773] = 12'b111111111111;
assign CPM[5774] = 12'b111111111111;
assign CPM[5775] = 12'b111111111111;
assign CPM[5776] = 12'b111111111111;
assign CPM[5777] = 12'b111111111111;
assign CPM[5778] = 12'b111111111111;
assign CPM[5779] = 12'b111111111111;
assign CPM[5780] = 12'b111111111111;
assign CPM[5781] = 12'b111111111111;
assign CPM[5782] = 12'b111111111111;
assign CPM[5783] = 12'b111111111111;
assign CPM[5784] = 12'b111111111111;
assign CPM[5785] = 12'b111111111111;
assign CPM[5786] = 12'b111111111111;
assign CPM[5787] = 12'b111111111111;
assign CPM[5788] = 12'b111111111111;
assign CPM[5789] = 12'b111111111111;
assign CPM[5790] = 12'b111111111111;
assign CPM[5791] = 12'b111111111111;
assign CPM[5792] = 12'b111111111111;
assign CPM[5793] = 12'b111111111111;
assign CPM[5794] = 12'b111111111111;
assign CPM[5795] = 12'b111111111111;
assign CPM[5796] = 12'b111111111111;
assign CPM[5797] = 12'b111111111111;
assign CPM[5798] = 12'b111111111111;
assign CPM[5799] = 12'b111111111111;
assign CPM[5800] = 12'b111111111111;
assign CPM[5801] = 12'b000000000000;
assign CPM[5802] = 12'b000000000000;
assign CPM[5803] = 12'b000000000000;
assign CPM[5804] = 12'b000000000000;
assign CPM[5805] = 12'b111111111111;
assign CPM[5806] = 12'b111111111111;
assign CPM[5807] = 12'b111111111111;
assign CPM[5808] = 12'b111111111111;
assign CPM[5809] = 12'b111111111111;
assign CPM[5810] = 12'b111111111111;
assign CPM[5811] = 12'b111111111111;
assign CPM[5812] = 12'b111111111111;
assign CPM[5813] = 12'b111111111111;
assign CPM[5814] = 12'b111111111111;
assign CPM[5815] = 12'b111111111111;
assign CPM[5816] = 12'b111111111111;
assign CPM[5817] = 12'b111111111111;
assign CPM[5818] = 12'b111111111111;
assign CPM[5819] = 12'b111111111111;
assign CPM[5820] = 12'b111111111111;
assign CPM[5821] = 12'b111111111111;
assign CPM[5822] = 12'b111111111111;
assign CPM[5823] = 12'b111111111111;
assign CPM[5824] = 12'b111111111111;
assign CPM[5825] = 12'b111111111111;
assign CPM[5826] = 12'b111111111111;
assign CPM[5827] = 12'b111111111111;
assign CPM[5828] = 12'b111111111111;
assign CPM[5829] = 12'b111111111111;
assign CPM[5830] = 12'b111111111111;
assign CPM[5831] = 12'b111111111111;
assign CPM[5832] = 12'b111111111111;
assign CPM[5833] = 12'b000000000000;
assign CPM[5834] = 12'b000000000000;
assign CPM[5835] = 12'b000000000000;
assign CPM[5836] = 12'b000000000000;
assign CPM[5837] = 12'b111111111111;
assign CPM[5838] = 12'b111111111111;
assign CPM[5839] = 12'b111111111111;
assign CPM[5840] = 12'b111111111111;
assign CPM[5841] = 12'b111111111111;
assign CPM[5842] = 12'b111111111111;
assign CPM[5843] = 12'b111111111111;
assign CPM[5844] = 12'b111111111111;
assign CPM[5845] = 12'b111111111111;
assign CPM[5846] = 12'b111111111111;
assign CPM[5847] = 12'b111111111111;
assign CPM[5848] = 12'b111111111111;
assign CPM[5849] = 12'b111111111111;
assign CPM[5850] = 12'b111111111111;
assign CPM[5851] = 12'b111111111111;
assign CPM[5852] = 12'b111111111111;
assign CPM[5853] = 12'b111111111111;
assign CPM[5854] = 12'b111111111111;
assign CPM[5855] = 12'b111111111111;
assign CPM[5856] = 12'b111111111111;
assign CPM[5857] = 12'b111111111111;
assign CPM[5858] = 12'b111111111111;
assign CPM[5859] = 12'b111111111111;
assign CPM[5860] = 12'b111111111111;
assign CPM[5861] = 12'b111111111111;
assign CPM[5862] = 12'b000000000000;
assign CPM[5863] = 12'b000000000000;
assign CPM[5864] = 12'b000000000000;
assign CPM[5865] = 12'b000000000000;
assign CPM[5866] = 12'b000000000000;
assign CPM[5867] = 12'b000000000000;
assign CPM[5868] = 12'b000000000000;
assign CPM[5869] = 12'b000000000000;
assign CPM[5870] = 12'b000000000000;
assign CPM[5871] = 12'b000000000000;
assign CPM[5872] = 12'b000000000000;
assign CPM[5873] = 12'b000000000000;
assign CPM[5874] = 12'b000000000000;
assign CPM[5875] = 12'b000000000000;
assign CPM[5876] = 12'b000000000000;
assign CPM[5877] = 12'b000000000000;
assign CPM[5878] = 12'b000000000000;
assign CPM[5879] = 12'b000000000000;
assign CPM[5880] = 12'b000000000000;
assign CPM[5881] = 12'b111111111111;
assign CPM[5882] = 12'b111111111111;
assign CPM[5883] = 12'b111111111111;
assign CPM[5884] = 12'b111111111111;
assign CPM[5885] = 12'b111111111111;
assign CPM[5886] = 12'b111111111111;
assign CPM[5887] = 12'b111111111111;
assign CPM[5888] = 12'b111111111111;
assign CPM[5889] = 12'b111111111111;
assign CPM[5890] = 12'b111111111111;
assign CPM[5891] = 12'b111111111111;
assign CPM[5892] = 12'b111111111111;
assign CPM[5893] = 12'b111111111111;
assign CPM[5894] = 12'b000000000000;
assign CPM[5895] = 12'b000000000000;
assign CPM[5896] = 12'b000000000000;
assign CPM[5897] = 12'b000000000000;
assign CPM[5898] = 12'b000000000000;
assign CPM[5899] = 12'b000000000000;
assign CPM[5900] = 12'b000000000000;
assign CPM[5901] = 12'b000000000000;
assign CPM[5902] = 12'b000000000000;
assign CPM[5903] = 12'b000000000000;
assign CPM[5904] = 12'b000000000000;
assign CPM[5905] = 12'b000000000000;
assign CPM[5906] = 12'b000000000000;
assign CPM[5907] = 12'b000000000000;
assign CPM[5908] = 12'b000000000000;
assign CPM[5909] = 12'b000000000000;
assign CPM[5910] = 12'b000000000000;
assign CPM[5911] = 12'b000000000000;
assign CPM[5912] = 12'b000000000000;
assign CPM[5913] = 12'b111111111111;
assign CPM[5914] = 12'b111111111111;
assign CPM[5915] = 12'b111111111111;
assign CPM[5916] = 12'b111111111111;
assign CPM[5917] = 12'b111111111111;
assign CPM[5918] = 12'b111111111111;
assign CPM[5919] = 12'b111111111111;
assign CPM[5920] = 12'b111111111111;
assign CPM[5921] = 12'b111111111111;
assign CPM[5922] = 12'b111111111111;
assign CPM[5923] = 12'b111111111111;
assign CPM[5924] = 12'b111111111111;
assign CPM[5925] = 12'b111111111111;
assign CPM[5926] = 12'b000000000000;
assign CPM[5927] = 12'b000000000000;
assign CPM[5928] = 12'b000000000000;
assign CPM[5929] = 12'b000000000000;
assign CPM[5930] = 12'b000000000000;
assign CPM[5931] = 12'b000000000000;
assign CPM[5932] = 12'b000000000000;
assign CPM[5933] = 12'b000000000000;
assign CPM[5934] = 12'b000000000000;
assign CPM[5935] = 12'b000000000000;
assign CPM[5936] = 12'b000000000000;
assign CPM[5937] = 12'b000000000000;
assign CPM[5938] = 12'b000000000000;
assign CPM[5939] = 12'b000000000000;
assign CPM[5940] = 12'b000000000000;
assign CPM[5941] = 12'b000000000000;
assign CPM[5942] = 12'b000000000000;
assign CPM[5943] = 12'b000000000000;
assign CPM[5944] = 12'b000000000000;
assign CPM[5945] = 12'b111111111111;
assign CPM[5946] = 12'b111111111111;
assign CPM[5947] = 12'b111111111111;
assign CPM[5948] = 12'b111111111111;
assign CPM[5949] = 12'b111111111111;
assign CPM[5950] = 12'b111111111111;
assign CPM[5951] = 12'b111111111111;
assign CPM[5952] = 12'b111111111111;
assign CPM[5953] = 12'b111111111111;
assign CPM[5954] = 12'b111111111111;
assign CPM[5955] = 12'b111111111111;
assign CPM[5956] = 12'b111111111111;
assign CPM[5957] = 12'b111111111111;
assign CPM[5958] = 12'b000000000000;
assign CPM[5959] = 12'b000000000000;
assign CPM[5960] = 12'b000000000000;
assign CPM[5961] = 12'b000000000000;
assign CPM[5962] = 12'b000000000000;
assign CPM[5963] = 12'b000000000000;
assign CPM[5964] = 12'b000000000000;
assign CPM[5965] = 12'b000000000000;
assign CPM[5966] = 12'b000000000000;
assign CPM[5967] = 12'b000000000000;
assign CPM[5968] = 12'b000000000000;
assign CPM[5969] = 12'b000000000000;
assign CPM[5970] = 12'b000000000000;
assign CPM[5971] = 12'b000000000000;
assign CPM[5972] = 12'b000000000000;
assign CPM[5973] = 12'b000000000000;
assign CPM[5974] = 12'b000000000000;
assign CPM[5975] = 12'b000000000000;
assign CPM[5976] = 12'b000000000000;
assign CPM[5977] = 12'b111111111111;
assign CPM[5978] = 12'b111111111111;
assign CPM[5979] = 12'b111111111111;
assign CPM[5980] = 12'b111111111111;
assign CPM[5981] = 12'b111111111111;
assign CPM[5982] = 12'b111111111111;
assign CPM[5983] = 12'b111111111111;
assign CPM[5984] = 12'b111111111111;
assign CPM[5985] = 12'b111111111111;
assign CPM[5986] = 12'b111111111111;
assign CPM[5987] = 12'b111111111111;
assign CPM[5988] = 12'b111111111111;
assign CPM[5989] = 12'b111111111111;
assign CPM[5990] = 12'b111111111111;
assign CPM[5991] = 12'b111111111111;
assign CPM[5992] = 12'b111111111111;
assign CPM[5993] = 12'b111111111111;
assign CPM[5994] = 12'b111111111111;
assign CPM[5995] = 12'b111111111111;
assign CPM[5996] = 12'b111111111111;
assign CPM[5997] = 12'b111111111111;
assign CPM[5998] = 12'b111111111111;
assign CPM[5999] = 12'b111111111111;
assign CPM[6000] = 12'b111111111111;
assign CPM[6001] = 12'b111111111111;
assign CPM[6002] = 12'b111111111111;
assign CPM[6003] = 12'b111111111111;
assign CPM[6004] = 12'b111111111111;
assign CPM[6005] = 12'b111111111111;
assign CPM[6006] = 12'b111111111111;
assign CPM[6007] = 12'b111111111111;
assign CPM[6008] = 12'b111111111111;
assign CPM[6009] = 12'b111111111111;
assign CPM[6010] = 12'b111111111111;
assign CPM[6011] = 12'b111111111111;
assign CPM[6012] = 12'b111111111111;
assign CPM[6013] = 12'b111111111111;
assign CPM[6014] = 12'b111111111111;
assign CPM[6015] = 12'b111111111111;
assign CPM[6016] = 12'b111111111111;
assign CPM[6017] = 12'b111111111111;
assign CPM[6018] = 12'b111111111111;
assign CPM[6019] = 12'b111111111111;
assign CPM[6020] = 12'b111111111111;
assign CPM[6021] = 12'b111111111111;
assign CPM[6022] = 12'b111111111111;
assign CPM[6023] = 12'b111111111111;
assign CPM[6024] = 12'b111111111111;
assign CPM[6025] = 12'b111111111111;
assign CPM[6026] = 12'b111111111111;
assign CPM[6027] = 12'b111111111111;
assign CPM[6028] = 12'b111111111111;
assign CPM[6029] = 12'b111111111111;
assign CPM[6030] = 12'b111111111111;
assign CPM[6031] = 12'b111111111111;
assign CPM[6032] = 12'b111111111111;
assign CPM[6033] = 12'b111111111111;
assign CPM[6034] = 12'b111111111111;
assign CPM[6035] = 12'b111111111111;
assign CPM[6036] = 12'b111111111111;
assign CPM[6037] = 12'b111111111111;
assign CPM[6038] = 12'b111111111111;
assign CPM[6039] = 12'b111111111111;
assign CPM[6040] = 12'b111111111111;
assign CPM[6041] = 12'b111111111111;
assign CPM[6042] = 12'b111111111111;
assign CPM[6043] = 12'b111111111111;
assign CPM[6044] = 12'b111111111111;
assign CPM[6045] = 12'b111111111111;
assign CPM[6046] = 12'b111111111111;
assign CPM[6047] = 12'b111111111111;
assign CPM[6048] = 12'b111111111111;
assign CPM[6049] = 12'b111111111111;
assign CPM[6050] = 12'b111111111111;
assign CPM[6051] = 12'b111111111111;
assign CPM[6052] = 12'b111111111111;
assign CPM[6053] = 12'b111111111111;
assign CPM[6054] = 12'b111111111111;
assign CPM[6055] = 12'b111111111111;
assign CPM[6056] = 12'b111111111111;
assign CPM[6057] = 12'b111111111111;
assign CPM[6058] = 12'b111111111111;
assign CPM[6059] = 12'b111111111111;
assign CPM[6060] = 12'b111111111111;
assign CPM[6061] = 12'b111111111111;
assign CPM[6062] = 12'b111111111111;
assign CPM[6063] = 12'b111111111111;
assign CPM[6064] = 12'b111111111111;
assign CPM[6065] = 12'b111111111111;
assign CPM[6066] = 12'b111111111111;
assign CPM[6067] = 12'b111111111111;
assign CPM[6068] = 12'b111111111111;
assign CPM[6069] = 12'b111111111111;
assign CPM[6070] = 12'b111111111111;
assign CPM[6071] = 12'b111111111111;
assign CPM[6072] = 12'b111111111111;
assign CPM[6073] = 12'b111111111111;
assign CPM[6074] = 12'b111111111111;
assign CPM[6075] = 12'b111111111111;
assign CPM[6076] = 12'b111111111111;
assign CPM[6077] = 12'b111111111111;
assign CPM[6078] = 12'b111111111111;
assign CPM[6079] = 12'b111111111111;
assign CPM[6080] = 12'b111111111111;
assign CPM[6081] = 12'b111111111111;
assign CPM[6082] = 12'b111111111111;
assign CPM[6083] = 12'b111111111111;
assign CPM[6084] = 12'b111111111111;
assign CPM[6085] = 12'b111111111111;
assign CPM[6086] = 12'b111111111111;
assign CPM[6087] = 12'b111111111111;
assign CPM[6088] = 12'b111111111111;
assign CPM[6089] = 12'b111111111111;
assign CPM[6090] = 12'b111111111111;
assign CPM[6091] = 12'b111111111111;
assign CPM[6092] = 12'b111111111111;
assign CPM[6093] = 12'b111111111111;
assign CPM[6094] = 12'b111111111111;
assign CPM[6095] = 12'b111111111111;
assign CPM[6096] = 12'b111111111111;
assign CPM[6097] = 12'b111111111111;
assign CPM[6098] = 12'b111111111111;
assign CPM[6099] = 12'b111111111111;
assign CPM[6100] = 12'b111111111111;
assign CPM[6101] = 12'b111111111111;
assign CPM[6102] = 12'b111111111111;
assign CPM[6103] = 12'b111111111111;
assign CPM[6104] = 12'b111111111111;
assign CPM[6105] = 12'b111111111111;
assign CPM[6106] = 12'b111111111111;
assign CPM[6107] = 12'b111111111111;
assign CPM[6108] = 12'b111111111111;
assign CPM[6109] = 12'b111111111111;
assign CPM[6110] = 12'b111111111111;
assign CPM[6111] = 12'b111111111111;
assign CPM[6112] = 12'b111111111111;
assign CPM[6113] = 12'b111111111111;
assign CPM[6114] = 12'b111111111111;
assign CPM[6115] = 12'b111111111111;
assign CPM[6116] = 12'b111111111111;
assign CPM[6117] = 12'b111111111111;
assign CPM[6118] = 12'b111111111111;
assign CPM[6119] = 12'b111111111111;
assign CPM[6120] = 12'b111111111111;
assign CPM[6121] = 12'b111111111111;
assign CPM[6122] = 12'b111111111111;
assign CPM[6123] = 12'b111111111111;
assign CPM[6124] = 12'b111111111111;
assign CPM[6125] = 12'b111111111111;
assign CPM[6126] = 12'b111111111111;
assign CPM[6127] = 12'b111111111111;
assign CPM[6128] = 12'b111111111111;
assign CPM[6129] = 12'b111111111111;
assign CPM[6130] = 12'b111111111111;
assign CPM[6131] = 12'b111111111111;
assign CPM[6132] = 12'b111111111111;
assign CPM[6133] = 12'b111111111111;
assign CPM[6134] = 12'b111111111111;
assign CPM[6135] = 12'b111111111111;
assign CPM[6136] = 12'b111111111111;
assign CPM[6137] = 12'b111111111111;
assign CPM[6138] = 12'b111111111111;
assign CPM[6139] = 12'b111111111111;
assign CPM[6140] = 12'b111111111111;
assign CPM[6141] = 12'b111111111111;
assign CPM[6142] = 12'b111111111111;
assign CPM[6143] = 12'b111111111111;
assign CPM[6144] = 12'b111111111111;
assign CPM[6145] = 12'b111111111111;
assign CPM[6146] = 12'b111111111111;
assign CPM[6147] = 12'b111111111111;
assign CPM[6148] = 12'b111111111111;
assign CPM[6149] = 12'b111111111111;
assign CPM[6150] = 12'b111111111111;
assign CPM[6151] = 12'b111111111111;
assign CPM[6152] = 12'b111111111111;
assign CPM[6153] = 12'b111111111111;
assign CPM[6154] = 12'b111111111111;
assign CPM[6155] = 12'b111111111111;
assign CPM[6156] = 12'b111111111111;
assign CPM[6157] = 12'b111111111111;
assign CPM[6158] = 12'b111111111111;
assign CPM[6159] = 12'b111111111111;
assign CPM[6160] = 12'b111111111111;
assign CPM[6161] = 12'b111111111111;
assign CPM[6162] = 12'b111111111111;
assign CPM[6163] = 12'b111111111111;
assign CPM[6164] = 12'b111111111111;
assign CPM[6165] = 12'b111111111111;
assign CPM[6166] = 12'b111111111111;
assign CPM[6167] = 12'b111111111111;
assign CPM[6168] = 12'b111111111111;
assign CPM[6169] = 12'b111111111111;
assign CPM[6170] = 12'b111111111111;
assign CPM[6171] = 12'b111111111111;
assign CPM[6172] = 12'b111111111111;
assign CPM[6173] = 12'b111111111111;
assign CPM[6174] = 12'b111111111111;
assign CPM[6175] = 12'b111111111111;
assign CPM[6176] = 12'b111111111111;
assign CPM[6177] = 12'b111111111111;
assign CPM[6178] = 12'b111111111111;
assign CPM[6179] = 12'b111111111111;
assign CPM[6180] = 12'b111111111111;
assign CPM[6181] = 12'b111111111111;
assign CPM[6182] = 12'b111111111111;
assign CPM[6183] = 12'b111111111111;
assign CPM[6184] = 12'b111111111111;
assign CPM[6185] = 12'b111111111111;
assign CPM[6186] = 12'b111111111111;
assign CPM[6187] = 12'b111111111111;
assign CPM[6188] = 12'b111111111111;
assign CPM[6189] = 12'b111111111111;
assign CPM[6190] = 12'b111111111111;
assign CPM[6191] = 12'b111111111111;
assign CPM[6192] = 12'b111111111111;
assign CPM[6193] = 12'b111111111111;
assign CPM[6194] = 12'b111111111111;
assign CPM[6195] = 12'b111111111111;
assign CPM[6196] = 12'b111111111111;
assign CPM[6197] = 12'b111111111111;
assign CPM[6198] = 12'b111111111111;
assign CPM[6199] = 12'b111111111111;
assign CPM[6200] = 12'b111111111111;
assign CPM[6201] = 12'b111111111111;
assign CPM[6202] = 12'b111111111111;
assign CPM[6203] = 12'b111111111111;
assign CPM[6204] = 12'b111111111111;
assign CPM[6205] = 12'b111111111111;
assign CPM[6206] = 12'b111111111111;
assign CPM[6207] = 12'b111111111111;
assign CPM[6208] = 12'b111111111111;
assign CPM[6209] = 12'b111111111111;
assign CPM[6210] = 12'b111111111111;
assign CPM[6211] = 12'b111111111111;
assign CPM[6212] = 12'b111111111111;
assign CPM[6213] = 12'b111111111111;
assign CPM[6214] = 12'b111111111111;
assign CPM[6215] = 12'b111111111111;
assign CPM[6216] = 12'b111111111111;
assign CPM[6217] = 12'b111111111111;
assign CPM[6218] = 12'b111111111111;
assign CPM[6219] = 12'b000000000000;
assign CPM[6220] = 12'b000000000000;
assign CPM[6221] = 12'b000000000000;
assign CPM[6222] = 12'b000000000000;
assign CPM[6223] = 12'b000000000000;
assign CPM[6224] = 12'b000000000000;
assign CPM[6225] = 12'b000000000000;
assign CPM[6226] = 12'b000000000000;
assign CPM[6227] = 12'b000000000000;
assign CPM[6228] = 12'b000000000000;
assign CPM[6229] = 12'b111111111111;
assign CPM[6230] = 12'b111111111111;
assign CPM[6231] = 12'b111111111111;
assign CPM[6232] = 12'b111111111111;
assign CPM[6233] = 12'b111111111111;
assign CPM[6234] = 12'b111111111111;
assign CPM[6235] = 12'b111111111111;
assign CPM[6236] = 12'b111111111111;
assign CPM[6237] = 12'b111111111111;
assign CPM[6238] = 12'b111111111111;
assign CPM[6239] = 12'b111111111111;
assign CPM[6240] = 12'b111111111111;
assign CPM[6241] = 12'b111111111111;
assign CPM[6242] = 12'b111111111111;
assign CPM[6243] = 12'b111111111111;
assign CPM[6244] = 12'b111111111111;
assign CPM[6245] = 12'b111111111111;
assign CPM[6246] = 12'b111111111111;
assign CPM[6247] = 12'b111111111111;
assign CPM[6248] = 12'b111111111111;
assign CPM[6249] = 12'b111111111111;
assign CPM[6250] = 12'b111111111111;
assign CPM[6251] = 12'b000000000000;
assign CPM[6252] = 12'b000000000000;
assign CPM[6253] = 12'b000000000000;
assign CPM[6254] = 12'b000000000000;
assign CPM[6255] = 12'b000000000000;
assign CPM[6256] = 12'b000000000000;
assign CPM[6257] = 12'b000000000000;
assign CPM[6258] = 12'b000000000000;
assign CPM[6259] = 12'b000000000000;
assign CPM[6260] = 12'b000000000000;
assign CPM[6261] = 12'b111111111111;
assign CPM[6262] = 12'b111111111111;
assign CPM[6263] = 12'b111111111111;
assign CPM[6264] = 12'b111111111111;
assign CPM[6265] = 12'b111111111111;
assign CPM[6266] = 12'b111111111111;
assign CPM[6267] = 12'b111111111111;
assign CPM[6268] = 12'b111111111111;
assign CPM[6269] = 12'b111111111111;
assign CPM[6270] = 12'b111111111111;
assign CPM[6271] = 12'b111111111111;
assign CPM[6272] = 12'b111111111111;
assign CPM[6273] = 12'b111111111111;
assign CPM[6274] = 12'b111111111111;
assign CPM[6275] = 12'b111111111111;
assign CPM[6276] = 12'b111111111111;
assign CPM[6277] = 12'b111111111111;
assign CPM[6278] = 12'b111111111111;
assign CPM[6279] = 12'b111111111111;
assign CPM[6280] = 12'b111111111111;
assign CPM[6281] = 12'b111111111111;
assign CPM[6282] = 12'b111111111111;
assign CPM[6283] = 12'b000000000000;
assign CPM[6284] = 12'b000000000000;
assign CPM[6285] = 12'b000000000000;
assign CPM[6286] = 12'b000000000000;
assign CPM[6287] = 12'b000000000000;
assign CPM[6288] = 12'b000000000000;
assign CPM[6289] = 12'b000000000000;
assign CPM[6290] = 12'b000000000000;
assign CPM[6291] = 12'b000000000000;
assign CPM[6292] = 12'b000000000000;
assign CPM[6293] = 12'b111111111111;
assign CPM[6294] = 12'b111111111111;
assign CPM[6295] = 12'b111111111111;
assign CPM[6296] = 12'b111111111111;
assign CPM[6297] = 12'b111111111111;
assign CPM[6298] = 12'b111111111111;
assign CPM[6299] = 12'b111111111111;
assign CPM[6300] = 12'b111111111111;
assign CPM[6301] = 12'b111111111111;
assign CPM[6302] = 12'b111111111111;
assign CPM[6303] = 12'b111111111111;
assign CPM[6304] = 12'b111111111111;
assign CPM[6305] = 12'b111111111111;
assign CPM[6306] = 12'b111111111111;
assign CPM[6307] = 12'b111111111111;
assign CPM[6308] = 12'b111111111111;
assign CPM[6309] = 12'b111111111111;
assign CPM[6310] = 12'b111111111111;
assign CPM[6311] = 12'b111111111111;
assign CPM[6312] = 12'b111111111111;
assign CPM[6313] = 12'b111111111111;
assign CPM[6314] = 12'b111111111111;
assign CPM[6315] = 12'b000000000000;
assign CPM[6316] = 12'b000000000000;
assign CPM[6317] = 12'b000000000000;
assign CPM[6318] = 12'b000000000000;
assign CPM[6319] = 12'b000000000000;
assign CPM[6320] = 12'b000000000000;
assign CPM[6321] = 12'b000000000000;
assign CPM[6322] = 12'b000000000000;
assign CPM[6323] = 12'b000000000000;
assign CPM[6324] = 12'b000000000000;
assign CPM[6325] = 12'b111111111111;
assign CPM[6326] = 12'b111111111111;
assign CPM[6327] = 12'b111111111111;
assign CPM[6328] = 12'b111111111111;
assign CPM[6329] = 12'b111111111111;
assign CPM[6330] = 12'b111111111111;
assign CPM[6331] = 12'b111111111111;
assign CPM[6332] = 12'b111111111111;
assign CPM[6333] = 12'b111111111111;
assign CPM[6334] = 12'b111111111111;
assign CPM[6335] = 12'b111111111111;
assign CPM[6336] = 12'b111111111111;
assign CPM[6337] = 12'b111111111111;
assign CPM[6338] = 12'b111111111111;
assign CPM[6339] = 12'b111111111111;
assign CPM[6340] = 12'b111111111111;
assign CPM[6341] = 12'b111111111111;
assign CPM[6342] = 12'b111111111111;
assign CPM[6343] = 12'b000000000000;
assign CPM[6344] = 12'b000000000000;
assign CPM[6345] = 12'b000000000000;
assign CPM[6346] = 12'b000000000000;
assign CPM[6347] = 12'b111111111111;
assign CPM[6348] = 12'b111111111111;
assign CPM[6349] = 12'b111111111111;
assign CPM[6350] = 12'b111111111111;
assign CPM[6351] = 12'b111111111111;
assign CPM[6352] = 12'b111111111111;
assign CPM[6353] = 12'b111111111111;
assign CPM[6354] = 12'b111111111111;
assign CPM[6355] = 12'b111111111111;
assign CPM[6356] = 12'b111111111111;
assign CPM[6357] = 12'b000000000000;
assign CPM[6358] = 12'b000000000000;
assign CPM[6359] = 12'b000000000000;
assign CPM[6360] = 12'b000000000000;
assign CPM[6361] = 12'b111111111111;
assign CPM[6362] = 12'b111111111111;
assign CPM[6363] = 12'b111111111111;
assign CPM[6364] = 12'b111111111111;
assign CPM[6365] = 12'b111111111111;
assign CPM[6366] = 12'b111111111111;
assign CPM[6367] = 12'b111111111111;
assign CPM[6368] = 12'b111111111111;
assign CPM[6369] = 12'b111111111111;
assign CPM[6370] = 12'b111111111111;
assign CPM[6371] = 12'b111111111111;
assign CPM[6372] = 12'b111111111111;
assign CPM[6373] = 12'b111111111111;
assign CPM[6374] = 12'b111111111111;
assign CPM[6375] = 12'b000000000000;
assign CPM[6376] = 12'b000000000000;
assign CPM[6377] = 12'b000000000000;
assign CPM[6378] = 12'b000000000000;
assign CPM[6379] = 12'b111111111111;
assign CPM[6380] = 12'b111111111111;
assign CPM[6381] = 12'b111111111111;
assign CPM[6382] = 12'b111111111111;
assign CPM[6383] = 12'b111111111111;
assign CPM[6384] = 12'b111111111111;
assign CPM[6385] = 12'b111111111111;
assign CPM[6386] = 12'b111111111111;
assign CPM[6387] = 12'b111111111111;
assign CPM[6388] = 12'b111111111111;
assign CPM[6389] = 12'b000000000000;
assign CPM[6390] = 12'b000000000000;
assign CPM[6391] = 12'b000000000000;
assign CPM[6392] = 12'b000000000000;
assign CPM[6393] = 12'b111111111111;
assign CPM[6394] = 12'b111111111111;
assign CPM[6395] = 12'b111111111111;
assign CPM[6396] = 12'b111111111111;
assign CPM[6397] = 12'b111111111111;
assign CPM[6398] = 12'b111111111111;
assign CPM[6399] = 12'b111111111111;
assign CPM[6400] = 12'b111111111111;
assign CPM[6401] = 12'b111111111111;
assign CPM[6402] = 12'b111111111111;
assign CPM[6403] = 12'b111111111111;
assign CPM[6404] = 12'b111111111111;
assign CPM[6405] = 12'b111111111111;
assign CPM[6406] = 12'b111111111111;
assign CPM[6407] = 12'b000000000000;
assign CPM[6408] = 12'b000000000000;
assign CPM[6409] = 12'b000000000000;
assign CPM[6410] = 12'b000000000000;
assign CPM[6411] = 12'b111111111111;
assign CPM[6412] = 12'b111111111111;
assign CPM[6413] = 12'b111111111111;
assign CPM[6414] = 12'b111111111111;
assign CPM[6415] = 12'b111111111111;
assign CPM[6416] = 12'b111111111111;
assign CPM[6417] = 12'b111111111111;
assign CPM[6418] = 12'b111111111111;
assign CPM[6419] = 12'b111111111111;
assign CPM[6420] = 12'b111111111111;
assign CPM[6421] = 12'b000000000000;
assign CPM[6422] = 12'b000000000000;
assign CPM[6423] = 12'b000000000000;
assign CPM[6424] = 12'b000000000000;
assign CPM[6425] = 12'b111111111111;
assign CPM[6426] = 12'b111111111111;
assign CPM[6427] = 12'b111111111111;
assign CPM[6428] = 12'b111111111111;
assign CPM[6429] = 12'b111111111111;
assign CPM[6430] = 12'b111111111111;
assign CPM[6431] = 12'b111111111111;
assign CPM[6432] = 12'b111111111111;
assign CPM[6433] = 12'b111111111111;
assign CPM[6434] = 12'b111111111111;
assign CPM[6435] = 12'b111111111111;
assign CPM[6436] = 12'b111111111111;
assign CPM[6437] = 12'b111111111111;
assign CPM[6438] = 12'b111111111111;
assign CPM[6439] = 12'b000000000000;
assign CPM[6440] = 12'b000000000000;
assign CPM[6441] = 12'b000000000000;
assign CPM[6442] = 12'b000000000000;
assign CPM[6443] = 12'b111111111111;
assign CPM[6444] = 12'b111111111111;
assign CPM[6445] = 12'b111111111111;
assign CPM[6446] = 12'b111111111111;
assign CPM[6447] = 12'b111111111111;
assign CPM[6448] = 12'b111111111111;
assign CPM[6449] = 12'b111111111111;
assign CPM[6450] = 12'b111111111111;
assign CPM[6451] = 12'b111111111111;
assign CPM[6452] = 12'b111111111111;
assign CPM[6453] = 12'b000000000000;
assign CPM[6454] = 12'b000000000000;
assign CPM[6455] = 12'b000000000000;
assign CPM[6456] = 12'b000000000000;
assign CPM[6457] = 12'b111111111111;
assign CPM[6458] = 12'b111111111111;
assign CPM[6459] = 12'b111111111111;
assign CPM[6460] = 12'b111111111111;
assign CPM[6461] = 12'b111111111111;
assign CPM[6462] = 12'b111111111111;
assign CPM[6463] = 12'b111111111111;
assign CPM[6464] = 12'b111111111111;
assign CPM[6465] = 12'b111111111111;
assign CPM[6466] = 12'b111111111111;
assign CPM[6467] = 12'b111111111111;
assign CPM[6468] = 12'b111111111111;
assign CPM[6469] = 12'b111111111111;
assign CPM[6470] = 12'b111111111111;
assign CPM[6471] = 12'b111111111111;
assign CPM[6472] = 12'b111111111111;
assign CPM[6473] = 12'b111111111111;
assign CPM[6474] = 12'b111111111111;
assign CPM[6475] = 12'b111111111111;
assign CPM[6476] = 12'b111111111111;
assign CPM[6477] = 12'b111111111111;
assign CPM[6478] = 12'b111111111111;
assign CPM[6479] = 12'b111111111111;
assign CPM[6480] = 12'b111111111111;
assign CPM[6481] = 12'b111111111111;
assign CPM[6482] = 12'b111111111111;
assign CPM[6483] = 12'b111111111111;
assign CPM[6484] = 12'b111111111111;
assign CPM[6485] = 12'b000000000000;
assign CPM[6486] = 12'b000000000000;
assign CPM[6487] = 12'b000000000000;
assign CPM[6488] = 12'b000000000000;
assign CPM[6489] = 12'b111111111111;
assign CPM[6490] = 12'b111111111111;
assign CPM[6491] = 12'b111111111111;
assign CPM[6492] = 12'b111111111111;
assign CPM[6493] = 12'b111111111111;
assign CPM[6494] = 12'b111111111111;
assign CPM[6495] = 12'b111111111111;
assign CPM[6496] = 12'b111111111111;
assign CPM[6497] = 12'b111111111111;
assign CPM[6498] = 12'b111111111111;
assign CPM[6499] = 12'b111111111111;
assign CPM[6500] = 12'b111111111111;
assign CPM[6501] = 12'b111111111111;
assign CPM[6502] = 12'b111111111111;
assign CPM[6503] = 12'b111111111111;
assign CPM[6504] = 12'b111111111111;
assign CPM[6505] = 12'b111111111111;
assign CPM[6506] = 12'b111111111111;
assign CPM[6507] = 12'b111111111111;
assign CPM[6508] = 12'b111111111111;
assign CPM[6509] = 12'b111111111111;
assign CPM[6510] = 12'b111111111111;
assign CPM[6511] = 12'b111111111111;
assign CPM[6512] = 12'b111111111111;
assign CPM[6513] = 12'b111111111111;
assign CPM[6514] = 12'b111111111111;
assign CPM[6515] = 12'b111111111111;
assign CPM[6516] = 12'b111111111111;
assign CPM[6517] = 12'b000000000000;
assign CPM[6518] = 12'b000000000000;
assign CPM[6519] = 12'b000000000000;
assign CPM[6520] = 12'b000000000000;
assign CPM[6521] = 12'b111111111111;
assign CPM[6522] = 12'b111111111111;
assign CPM[6523] = 12'b111111111111;
assign CPM[6524] = 12'b111111111111;
assign CPM[6525] = 12'b111111111111;
assign CPM[6526] = 12'b111111111111;
assign CPM[6527] = 12'b111111111111;
assign CPM[6528] = 12'b111111111111;
assign CPM[6529] = 12'b111111111111;
assign CPM[6530] = 12'b111111111111;
assign CPM[6531] = 12'b111111111111;
assign CPM[6532] = 12'b111111111111;
assign CPM[6533] = 12'b111111111111;
assign CPM[6534] = 12'b111111111111;
assign CPM[6535] = 12'b111111111111;
assign CPM[6536] = 12'b111111111111;
assign CPM[6537] = 12'b111111111111;
assign CPM[6538] = 12'b111111111111;
assign CPM[6539] = 12'b111111111111;
assign CPM[6540] = 12'b111111111111;
assign CPM[6541] = 12'b111111111111;
assign CPM[6542] = 12'b111111111111;
assign CPM[6543] = 12'b111111111111;
assign CPM[6544] = 12'b111111111111;
assign CPM[6545] = 12'b111111111111;
assign CPM[6546] = 12'b111111111111;
assign CPM[6547] = 12'b111111111111;
assign CPM[6548] = 12'b111111111111;
assign CPM[6549] = 12'b000000000000;
assign CPM[6550] = 12'b000000000000;
assign CPM[6551] = 12'b000000000000;
assign CPM[6552] = 12'b000000000000;
assign CPM[6553] = 12'b111111111111;
assign CPM[6554] = 12'b111111111111;
assign CPM[6555] = 12'b111111111111;
assign CPM[6556] = 12'b111111111111;
assign CPM[6557] = 12'b111111111111;
assign CPM[6558] = 12'b111111111111;
assign CPM[6559] = 12'b111111111111;
assign CPM[6560] = 12'b111111111111;
assign CPM[6561] = 12'b111111111111;
assign CPM[6562] = 12'b111111111111;
assign CPM[6563] = 12'b111111111111;
assign CPM[6564] = 12'b111111111111;
assign CPM[6565] = 12'b111111111111;
assign CPM[6566] = 12'b111111111111;
assign CPM[6567] = 12'b111111111111;
assign CPM[6568] = 12'b111111111111;
assign CPM[6569] = 12'b111111111111;
assign CPM[6570] = 12'b111111111111;
assign CPM[6571] = 12'b111111111111;
assign CPM[6572] = 12'b111111111111;
assign CPM[6573] = 12'b111111111111;
assign CPM[6574] = 12'b111111111111;
assign CPM[6575] = 12'b000000000000;
assign CPM[6576] = 12'b000000000000;
assign CPM[6577] = 12'b000000000000;
assign CPM[6578] = 12'b000000000000;
assign CPM[6579] = 12'b000000000000;
assign CPM[6580] = 12'b000000000000;
assign CPM[6581] = 12'b111111111111;
assign CPM[6582] = 12'b111111111111;
assign CPM[6583] = 12'b111111111111;
assign CPM[6584] = 12'b111111111111;
assign CPM[6585] = 12'b111111111111;
assign CPM[6586] = 12'b111111111111;
assign CPM[6587] = 12'b111111111111;
assign CPM[6588] = 12'b111111111111;
assign CPM[6589] = 12'b111111111111;
assign CPM[6590] = 12'b111111111111;
assign CPM[6591] = 12'b111111111111;
assign CPM[6592] = 12'b111111111111;
assign CPM[6593] = 12'b111111111111;
assign CPM[6594] = 12'b111111111111;
assign CPM[6595] = 12'b111111111111;
assign CPM[6596] = 12'b111111111111;
assign CPM[6597] = 12'b111111111111;
assign CPM[6598] = 12'b111111111111;
assign CPM[6599] = 12'b111111111111;
assign CPM[6600] = 12'b111111111111;
assign CPM[6601] = 12'b111111111111;
assign CPM[6602] = 12'b111111111111;
assign CPM[6603] = 12'b111111111111;
assign CPM[6604] = 12'b111111111111;
assign CPM[6605] = 12'b111111111111;
assign CPM[6606] = 12'b111111111111;
assign CPM[6607] = 12'b000000000000;
assign CPM[6608] = 12'b000000000000;
assign CPM[6609] = 12'b000000000000;
assign CPM[6610] = 12'b000000000000;
assign CPM[6611] = 12'b000000000000;
assign CPM[6612] = 12'b000000000000;
assign CPM[6613] = 12'b111111111111;
assign CPM[6614] = 12'b111111111111;
assign CPM[6615] = 12'b111111111111;
assign CPM[6616] = 12'b111111111111;
assign CPM[6617] = 12'b111111111111;
assign CPM[6618] = 12'b111111111111;
assign CPM[6619] = 12'b111111111111;
assign CPM[6620] = 12'b111111111111;
assign CPM[6621] = 12'b111111111111;
assign CPM[6622] = 12'b111111111111;
assign CPM[6623] = 12'b111111111111;
assign CPM[6624] = 12'b111111111111;
assign CPM[6625] = 12'b111111111111;
assign CPM[6626] = 12'b111111111111;
assign CPM[6627] = 12'b111111111111;
assign CPM[6628] = 12'b111111111111;
assign CPM[6629] = 12'b111111111111;
assign CPM[6630] = 12'b111111111111;
assign CPM[6631] = 12'b111111111111;
assign CPM[6632] = 12'b111111111111;
assign CPM[6633] = 12'b111111111111;
assign CPM[6634] = 12'b111111111111;
assign CPM[6635] = 12'b111111111111;
assign CPM[6636] = 12'b111111111111;
assign CPM[6637] = 12'b111111111111;
assign CPM[6638] = 12'b111111111111;
assign CPM[6639] = 12'b000000000000;
assign CPM[6640] = 12'b000000000000;
assign CPM[6641] = 12'b000000000000;
assign CPM[6642] = 12'b000000000000;
assign CPM[6643] = 12'b000000000000;
assign CPM[6644] = 12'b000000000000;
assign CPM[6645] = 12'b111111111111;
assign CPM[6646] = 12'b111111111111;
assign CPM[6647] = 12'b111111111111;
assign CPM[6648] = 12'b111111111111;
assign CPM[6649] = 12'b111111111111;
assign CPM[6650] = 12'b111111111111;
assign CPM[6651] = 12'b111111111111;
assign CPM[6652] = 12'b111111111111;
assign CPM[6653] = 12'b111111111111;
assign CPM[6654] = 12'b111111111111;
assign CPM[6655] = 12'b111111111111;
assign CPM[6656] = 12'b111111111111;
assign CPM[6657] = 12'b111111111111;
assign CPM[6658] = 12'b111111111111;
assign CPM[6659] = 12'b111111111111;
assign CPM[6660] = 12'b111111111111;
assign CPM[6661] = 12'b111111111111;
assign CPM[6662] = 12'b111111111111;
assign CPM[6663] = 12'b111111111111;
assign CPM[6664] = 12'b111111111111;
assign CPM[6665] = 12'b111111111111;
assign CPM[6666] = 12'b111111111111;
assign CPM[6667] = 12'b111111111111;
assign CPM[6668] = 12'b111111111111;
assign CPM[6669] = 12'b111111111111;
assign CPM[6670] = 12'b111111111111;
assign CPM[6671] = 12'b000000000000;
assign CPM[6672] = 12'b000000000000;
assign CPM[6673] = 12'b000000000000;
assign CPM[6674] = 12'b000000000000;
assign CPM[6675] = 12'b000000000000;
assign CPM[6676] = 12'b000000000000;
assign CPM[6677] = 12'b111111111111;
assign CPM[6678] = 12'b111111111111;
assign CPM[6679] = 12'b111111111111;
assign CPM[6680] = 12'b111111111111;
assign CPM[6681] = 12'b111111111111;
assign CPM[6682] = 12'b111111111111;
assign CPM[6683] = 12'b111111111111;
assign CPM[6684] = 12'b111111111111;
assign CPM[6685] = 12'b111111111111;
assign CPM[6686] = 12'b111111111111;
assign CPM[6687] = 12'b111111111111;
assign CPM[6688] = 12'b111111111111;
assign CPM[6689] = 12'b111111111111;
assign CPM[6690] = 12'b111111111111;
assign CPM[6691] = 12'b111111111111;
assign CPM[6692] = 12'b111111111111;
assign CPM[6693] = 12'b111111111111;
assign CPM[6694] = 12'b111111111111;
assign CPM[6695] = 12'b111111111111;
assign CPM[6696] = 12'b111111111111;
assign CPM[6697] = 12'b111111111111;
assign CPM[6698] = 12'b111111111111;
assign CPM[6699] = 12'b111111111111;
assign CPM[6700] = 12'b111111111111;
assign CPM[6701] = 12'b111111111111;
assign CPM[6702] = 12'b111111111111;
assign CPM[6703] = 12'b111111111111;
assign CPM[6704] = 12'b111111111111;
assign CPM[6705] = 12'b111111111111;
assign CPM[6706] = 12'b111111111111;
assign CPM[6707] = 12'b111111111111;
assign CPM[6708] = 12'b111111111111;
assign CPM[6709] = 12'b000000000000;
assign CPM[6710] = 12'b000000000000;
assign CPM[6711] = 12'b000000000000;
assign CPM[6712] = 12'b000000000000;
assign CPM[6713] = 12'b111111111111;
assign CPM[6714] = 12'b111111111111;
assign CPM[6715] = 12'b111111111111;
assign CPM[6716] = 12'b111111111111;
assign CPM[6717] = 12'b111111111111;
assign CPM[6718] = 12'b111111111111;
assign CPM[6719] = 12'b111111111111;
assign CPM[6720] = 12'b111111111111;
assign CPM[6721] = 12'b111111111111;
assign CPM[6722] = 12'b111111111111;
assign CPM[6723] = 12'b111111111111;
assign CPM[6724] = 12'b111111111111;
assign CPM[6725] = 12'b111111111111;
assign CPM[6726] = 12'b111111111111;
assign CPM[6727] = 12'b111111111111;
assign CPM[6728] = 12'b111111111111;
assign CPM[6729] = 12'b111111111111;
assign CPM[6730] = 12'b111111111111;
assign CPM[6731] = 12'b111111111111;
assign CPM[6732] = 12'b111111111111;
assign CPM[6733] = 12'b111111111111;
assign CPM[6734] = 12'b111111111111;
assign CPM[6735] = 12'b111111111111;
assign CPM[6736] = 12'b111111111111;
assign CPM[6737] = 12'b111111111111;
assign CPM[6738] = 12'b111111111111;
assign CPM[6739] = 12'b111111111111;
assign CPM[6740] = 12'b111111111111;
assign CPM[6741] = 12'b000000000000;
assign CPM[6742] = 12'b000000000000;
assign CPM[6743] = 12'b000000000000;
assign CPM[6744] = 12'b000000000000;
assign CPM[6745] = 12'b111111111111;
assign CPM[6746] = 12'b111111111111;
assign CPM[6747] = 12'b111111111111;
assign CPM[6748] = 12'b111111111111;
assign CPM[6749] = 12'b111111111111;
assign CPM[6750] = 12'b111111111111;
assign CPM[6751] = 12'b111111111111;
assign CPM[6752] = 12'b111111111111;
assign CPM[6753] = 12'b111111111111;
assign CPM[6754] = 12'b111111111111;
assign CPM[6755] = 12'b111111111111;
assign CPM[6756] = 12'b111111111111;
assign CPM[6757] = 12'b111111111111;
assign CPM[6758] = 12'b111111111111;
assign CPM[6759] = 12'b111111111111;
assign CPM[6760] = 12'b111111111111;
assign CPM[6761] = 12'b111111111111;
assign CPM[6762] = 12'b111111111111;
assign CPM[6763] = 12'b111111111111;
assign CPM[6764] = 12'b111111111111;
assign CPM[6765] = 12'b111111111111;
assign CPM[6766] = 12'b111111111111;
assign CPM[6767] = 12'b111111111111;
assign CPM[6768] = 12'b111111111111;
assign CPM[6769] = 12'b111111111111;
assign CPM[6770] = 12'b111111111111;
assign CPM[6771] = 12'b111111111111;
assign CPM[6772] = 12'b111111111111;
assign CPM[6773] = 12'b000000000000;
assign CPM[6774] = 12'b000000000000;
assign CPM[6775] = 12'b000000000000;
assign CPM[6776] = 12'b000000000000;
assign CPM[6777] = 12'b111111111111;
assign CPM[6778] = 12'b111111111111;
assign CPM[6779] = 12'b111111111111;
assign CPM[6780] = 12'b111111111111;
assign CPM[6781] = 12'b111111111111;
assign CPM[6782] = 12'b111111111111;
assign CPM[6783] = 12'b111111111111;
assign CPM[6784] = 12'b111111111111;
assign CPM[6785] = 12'b111111111111;
assign CPM[6786] = 12'b111111111111;
assign CPM[6787] = 12'b111111111111;
assign CPM[6788] = 12'b111111111111;
assign CPM[6789] = 12'b111111111111;
assign CPM[6790] = 12'b111111111111;
assign CPM[6791] = 12'b111111111111;
assign CPM[6792] = 12'b111111111111;
assign CPM[6793] = 12'b111111111111;
assign CPM[6794] = 12'b111111111111;
assign CPM[6795] = 12'b111111111111;
assign CPM[6796] = 12'b111111111111;
assign CPM[6797] = 12'b111111111111;
assign CPM[6798] = 12'b111111111111;
assign CPM[6799] = 12'b111111111111;
assign CPM[6800] = 12'b111111111111;
assign CPM[6801] = 12'b111111111111;
assign CPM[6802] = 12'b111111111111;
assign CPM[6803] = 12'b111111111111;
assign CPM[6804] = 12'b111111111111;
assign CPM[6805] = 12'b000000000000;
assign CPM[6806] = 12'b000000000000;
assign CPM[6807] = 12'b000000000000;
assign CPM[6808] = 12'b000000000000;
assign CPM[6809] = 12'b111111111111;
assign CPM[6810] = 12'b111111111111;
assign CPM[6811] = 12'b111111111111;
assign CPM[6812] = 12'b111111111111;
assign CPM[6813] = 12'b111111111111;
assign CPM[6814] = 12'b111111111111;
assign CPM[6815] = 12'b111111111111;
assign CPM[6816] = 12'b111111111111;
assign CPM[6817] = 12'b111111111111;
assign CPM[6818] = 12'b111111111111;
assign CPM[6819] = 12'b111111111111;
assign CPM[6820] = 12'b111111111111;
assign CPM[6821] = 12'b111111111111;
assign CPM[6822] = 12'b111111111111;
assign CPM[6823] = 12'b000000000000;
assign CPM[6824] = 12'b000000000000;
assign CPM[6825] = 12'b000000000000;
assign CPM[6826] = 12'b000000000000;
assign CPM[6827] = 12'b111111111111;
assign CPM[6828] = 12'b111111111111;
assign CPM[6829] = 12'b111111111111;
assign CPM[6830] = 12'b111111111111;
assign CPM[6831] = 12'b111111111111;
assign CPM[6832] = 12'b111111111111;
assign CPM[6833] = 12'b111111111111;
assign CPM[6834] = 12'b111111111111;
assign CPM[6835] = 12'b111111111111;
assign CPM[6836] = 12'b111111111111;
assign CPM[6837] = 12'b000000000000;
assign CPM[6838] = 12'b000000000000;
assign CPM[6839] = 12'b000000000000;
assign CPM[6840] = 12'b000000000000;
assign CPM[6841] = 12'b111111111111;
assign CPM[6842] = 12'b111111111111;
assign CPM[6843] = 12'b111111111111;
assign CPM[6844] = 12'b111111111111;
assign CPM[6845] = 12'b111111111111;
assign CPM[6846] = 12'b111111111111;
assign CPM[6847] = 12'b111111111111;
assign CPM[6848] = 12'b111111111111;
assign CPM[6849] = 12'b111111111111;
assign CPM[6850] = 12'b111111111111;
assign CPM[6851] = 12'b111111111111;
assign CPM[6852] = 12'b111111111111;
assign CPM[6853] = 12'b111111111111;
assign CPM[6854] = 12'b111111111111;
assign CPM[6855] = 12'b000000000000;
assign CPM[6856] = 12'b000000000000;
assign CPM[6857] = 12'b000000000000;
assign CPM[6858] = 12'b000000000000;
assign CPM[6859] = 12'b111111111111;
assign CPM[6860] = 12'b111111111111;
assign CPM[6861] = 12'b111111111111;
assign CPM[6862] = 12'b111111111111;
assign CPM[6863] = 12'b111111111111;
assign CPM[6864] = 12'b111111111111;
assign CPM[6865] = 12'b111111111111;
assign CPM[6866] = 12'b111111111111;
assign CPM[6867] = 12'b111111111111;
assign CPM[6868] = 12'b111111111111;
assign CPM[6869] = 12'b000000000000;
assign CPM[6870] = 12'b000000000000;
assign CPM[6871] = 12'b000000000000;
assign CPM[6872] = 12'b000000000000;
assign CPM[6873] = 12'b111111111111;
assign CPM[6874] = 12'b111111111111;
assign CPM[6875] = 12'b111111111111;
assign CPM[6876] = 12'b111111111111;
assign CPM[6877] = 12'b111111111111;
assign CPM[6878] = 12'b111111111111;
assign CPM[6879] = 12'b111111111111;
assign CPM[6880] = 12'b111111111111;
assign CPM[6881] = 12'b111111111111;
assign CPM[6882] = 12'b111111111111;
assign CPM[6883] = 12'b111111111111;
assign CPM[6884] = 12'b111111111111;
assign CPM[6885] = 12'b111111111111;
assign CPM[6886] = 12'b111111111111;
assign CPM[6887] = 12'b000000000000;
assign CPM[6888] = 12'b000000000000;
assign CPM[6889] = 12'b000000000000;
assign CPM[6890] = 12'b000000000000;
assign CPM[6891] = 12'b111111111111;
assign CPM[6892] = 12'b111111111111;
assign CPM[6893] = 12'b111111111111;
assign CPM[6894] = 12'b111111111111;
assign CPM[6895] = 12'b111111111111;
assign CPM[6896] = 12'b111111111111;
assign CPM[6897] = 12'b111111111111;
assign CPM[6898] = 12'b111111111111;
assign CPM[6899] = 12'b111111111111;
assign CPM[6900] = 12'b111111111111;
assign CPM[6901] = 12'b000000000000;
assign CPM[6902] = 12'b000000000000;
assign CPM[6903] = 12'b000000000000;
assign CPM[6904] = 12'b000000000000;
assign CPM[6905] = 12'b111111111111;
assign CPM[6906] = 12'b111111111111;
assign CPM[6907] = 12'b111111111111;
assign CPM[6908] = 12'b111111111111;
assign CPM[6909] = 12'b111111111111;
assign CPM[6910] = 12'b111111111111;
assign CPM[6911] = 12'b111111111111;
assign CPM[6912] = 12'b111111111111;
assign CPM[6913] = 12'b111111111111;
assign CPM[6914] = 12'b111111111111;
assign CPM[6915] = 12'b111111111111;
assign CPM[6916] = 12'b111111111111;
assign CPM[6917] = 12'b111111111111;
assign CPM[6918] = 12'b111111111111;
assign CPM[6919] = 12'b000000000000;
assign CPM[6920] = 12'b000000000000;
assign CPM[6921] = 12'b000000000000;
assign CPM[6922] = 12'b000000000000;
assign CPM[6923] = 12'b111111111111;
assign CPM[6924] = 12'b111111111111;
assign CPM[6925] = 12'b111111111111;
assign CPM[6926] = 12'b111111111111;
assign CPM[6927] = 12'b111111111111;
assign CPM[6928] = 12'b111111111111;
assign CPM[6929] = 12'b111111111111;
assign CPM[6930] = 12'b111111111111;
assign CPM[6931] = 12'b111111111111;
assign CPM[6932] = 12'b111111111111;
assign CPM[6933] = 12'b000000000000;
assign CPM[6934] = 12'b000000000000;
assign CPM[6935] = 12'b000000000000;
assign CPM[6936] = 12'b000000000000;
assign CPM[6937] = 12'b111111111111;
assign CPM[6938] = 12'b111111111111;
assign CPM[6939] = 12'b111111111111;
assign CPM[6940] = 12'b111111111111;
assign CPM[6941] = 12'b111111111111;
assign CPM[6942] = 12'b111111111111;
assign CPM[6943] = 12'b111111111111;
assign CPM[6944] = 12'b111111111111;
assign CPM[6945] = 12'b111111111111;
assign CPM[6946] = 12'b111111111111;
assign CPM[6947] = 12'b111111111111;
assign CPM[6948] = 12'b111111111111;
assign CPM[6949] = 12'b111111111111;
assign CPM[6950] = 12'b111111111111;
assign CPM[6951] = 12'b111111111111;
assign CPM[6952] = 12'b111111111111;
assign CPM[6953] = 12'b111111111111;
assign CPM[6954] = 12'b111111111111;
assign CPM[6955] = 12'b000000000000;
assign CPM[6956] = 12'b000000000000;
assign CPM[6957] = 12'b000000000000;
assign CPM[6958] = 12'b000000000000;
assign CPM[6959] = 12'b000000000000;
assign CPM[6960] = 12'b000000000000;
assign CPM[6961] = 12'b000000000000;
assign CPM[6962] = 12'b000000000000;
assign CPM[6963] = 12'b000000000000;
assign CPM[6964] = 12'b000000000000;
assign CPM[6965] = 12'b111111111111;
assign CPM[6966] = 12'b111111111111;
assign CPM[6967] = 12'b111111111111;
assign CPM[6968] = 12'b111111111111;
assign CPM[6969] = 12'b111111111111;
assign CPM[6970] = 12'b111111111111;
assign CPM[6971] = 12'b111111111111;
assign CPM[6972] = 12'b111111111111;
assign CPM[6973] = 12'b111111111111;
assign CPM[6974] = 12'b111111111111;
assign CPM[6975] = 12'b111111111111;
assign CPM[6976] = 12'b111111111111;
assign CPM[6977] = 12'b111111111111;
assign CPM[6978] = 12'b111111111111;
assign CPM[6979] = 12'b111111111111;
assign CPM[6980] = 12'b111111111111;
assign CPM[6981] = 12'b111111111111;
assign CPM[6982] = 12'b111111111111;
assign CPM[6983] = 12'b111111111111;
assign CPM[6984] = 12'b111111111111;
assign CPM[6985] = 12'b111111111111;
assign CPM[6986] = 12'b111111111111;
assign CPM[6987] = 12'b000000000000;
assign CPM[6988] = 12'b000000000000;
assign CPM[6989] = 12'b000000000000;
assign CPM[6990] = 12'b000000000000;
assign CPM[6991] = 12'b000000000000;
assign CPM[6992] = 12'b000000000000;
assign CPM[6993] = 12'b000000000000;
assign CPM[6994] = 12'b000000000000;
assign CPM[6995] = 12'b000000000000;
assign CPM[6996] = 12'b000000000000;
assign CPM[6997] = 12'b111111111111;
assign CPM[6998] = 12'b111111111111;
assign CPM[6999] = 12'b111111111111;
assign CPM[7000] = 12'b111111111111;
assign CPM[7001] = 12'b111111111111;
assign CPM[7002] = 12'b111111111111;
assign CPM[7003] = 12'b111111111111;
assign CPM[7004] = 12'b111111111111;
assign CPM[7005] = 12'b111111111111;
assign CPM[7006] = 12'b111111111111;
assign CPM[7007] = 12'b111111111111;
assign CPM[7008] = 12'b111111111111;
assign CPM[7009] = 12'b111111111111;
assign CPM[7010] = 12'b111111111111;
assign CPM[7011] = 12'b111111111111;
assign CPM[7012] = 12'b111111111111;
assign CPM[7013] = 12'b111111111111;
assign CPM[7014] = 12'b111111111111;
assign CPM[7015] = 12'b111111111111;
assign CPM[7016] = 12'b111111111111;
assign CPM[7017] = 12'b111111111111;
assign CPM[7018] = 12'b111111111111;
assign CPM[7019] = 12'b000000000000;
assign CPM[7020] = 12'b000000000000;
assign CPM[7021] = 12'b000000000000;
assign CPM[7022] = 12'b000000000000;
assign CPM[7023] = 12'b000000000000;
assign CPM[7024] = 12'b000000000000;
assign CPM[7025] = 12'b000000000000;
assign CPM[7026] = 12'b000000000000;
assign CPM[7027] = 12'b000000000000;
assign CPM[7028] = 12'b000000000000;
assign CPM[7029] = 12'b111111111111;
assign CPM[7030] = 12'b111111111111;
assign CPM[7031] = 12'b111111111111;
assign CPM[7032] = 12'b111111111111;
assign CPM[7033] = 12'b111111111111;
assign CPM[7034] = 12'b111111111111;
assign CPM[7035] = 12'b111111111111;
assign CPM[7036] = 12'b111111111111;
assign CPM[7037] = 12'b111111111111;
assign CPM[7038] = 12'b111111111111;
assign CPM[7039] = 12'b111111111111;
assign CPM[7040] = 12'b111111111111;
assign CPM[7041] = 12'b111111111111;
assign CPM[7042] = 12'b111111111111;
assign CPM[7043] = 12'b111111111111;
assign CPM[7044] = 12'b111111111111;
assign CPM[7045] = 12'b111111111111;
assign CPM[7046] = 12'b111111111111;
assign CPM[7047] = 12'b111111111111;
assign CPM[7048] = 12'b111111111111;
assign CPM[7049] = 12'b111111111111;
assign CPM[7050] = 12'b111111111111;
assign CPM[7051] = 12'b000000000000;
assign CPM[7052] = 12'b000000000000;
assign CPM[7053] = 12'b000000000000;
assign CPM[7054] = 12'b000000000000;
assign CPM[7055] = 12'b000000000000;
assign CPM[7056] = 12'b000000000000;
assign CPM[7057] = 12'b000000000000;
assign CPM[7058] = 12'b000000000000;
assign CPM[7059] = 12'b000000000000;
assign CPM[7060] = 12'b000000000000;
assign CPM[7061] = 12'b111111111111;
assign CPM[7062] = 12'b111111111111;
assign CPM[7063] = 12'b111111111111;
assign CPM[7064] = 12'b111111111111;
assign CPM[7065] = 12'b111111111111;
assign CPM[7066] = 12'b111111111111;
assign CPM[7067] = 12'b111111111111;
assign CPM[7068] = 12'b111111111111;
assign CPM[7069] = 12'b111111111111;
assign CPM[7070] = 12'b111111111111;
assign CPM[7071] = 12'b111111111111;
assign CPM[7072] = 12'b111111111111;
assign CPM[7073] = 12'b111111111111;
assign CPM[7074] = 12'b111111111111;
assign CPM[7075] = 12'b111111111111;
assign CPM[7076] = 12'b111111111111;
assign CPM[7077] = 12'b111111111111;
assign CPM[7078] = 12'b111111111111;
assign CPM[7079] = 12'b111111111111;
assign CPM[7080] = 12'b111111111111;
assign CPM[7081] = 12'b111111111111;
assign CPM[7082] = 12'b111111111111;
assign CPM[7083] = 12'b111111111111;
assign CPM[7084] = 12'b111111111111;
assign CPM[7085] = 12'b111111111111;
assign CPM[7086] = 12'b111111111111;
assign CPM[7087] = 12'b111111111111;
assign CPM[7088] = 12'b111111111111;
assign CPM[7089] = 12'b111111111111;
assign CPM[7090] = 12'b111111111111;
assign CPM[7091] = 12'b111111111111;
assign CPM[7092] = 12'b111111111111;
assign CPM[7093] = 12'b111111111111;
assign CPM[7094] = 12'b111111111111;
assign CPM[7095] = 12'b111111111111;
assign CPM[7096] = 12'b111111111111;
assign CPM[7097] = 12'b111111111111;
assign CPM[7098] = 12'b111111111111;
assign CPM[7099] = 12'b111111111111;
assign CPM[7100] = 12'b111111111111;
assign CPM[7101] = 12'b111111111111;
assign CPM[7102] = 12'b111111111111;
assign CPM[7103] = 12'b111111111111;
assign CPM[7104] = 12'b111111111111;
assign CPM[7105] = 12'b111111111111;
assign CPM[7106] = 12'b111111111111;
assign CPM[7107] = 12'b111111111111;
assign CPM[7108] = 12'b111111111111;
assign CPM[7109] = 12'b111111111111;
assign CPM[7110] = 12'b111111111111;
assign CPM[7111] = 12'b111111111111;
assign CPM[7112] = 12'b111111111111;
assign CPM[7113] = 12'b111111111111;
assign CPM[7114] = 12'b111111111111;
assign CPM[7115] = 12'b111111111111;
assign CPM[7116] = 12'b111111111111;
assign CPM[7117] = 12'b111111111111;
assign CPM[7118] = 12'b111111111111;
assign CPM[7119] = 12'b111111111111;
assign CPM[7120] = 12'b111111111111;
assign CPM[7121] = 12'b111111111111;
assign CPM[7122] = 12'b111111111111;
assign CPM[7123] = 12'b111111111111;
assign CPM[7124] = 12'b111111111111;
assign CPM[7125] = 12'b111111111111;
assign CPM[7126] = 12'b111111111111;
assign CPM[7127] = 12'b111111111111;
assign CPM[7128] = 12'b111111111111;
assign CPM[7129] = 12'b111111111111;
assign CPM[7130] = 12'b111111111111;
assign CPM[7131] = 12'b111111111111;
assign CPM[7132] = 12'b111111111111;
assign CPM[7133] = 12'b111111111111;
assign CPM[7134] = 12'b111111111111;
assign CPM[7135] = 12'b111111111111;
assign CPM[7136] = 12'b111111111111;
assign CPM[7137] = 12'b111111111111;
assign CPM[7138] = 12'b111111111111;
assign CPM[7139] = 12'b111111111111;
assign CPM[7140] = 12'b111111111111;
assign CPM[7141] = 12'b111111111111;
assign CPM[7142] = 12'b111111111111;
assign CPM[7143] = 12'b111111111111;
assign CPM[7144] = 12'b111111111111;
assign CPM[7145] = 12'b111111111111;
assign CPM[7146] = 12'b111111111111;
assign CPM[7147] = 12'b111111111111;
assign CPM[7148] = 12'b111111111111;
assign CPM[7149] = 12'b111111111111;
assign CPM[7150] = 12'b111111111111;
assign CPM[7151] = 12'b111111111111;
assign CPM[7152] = 12'b111111111111;
assign CPM[7153] = 12'b111111111111;
assign CPM[7154] = 12'b111111111111;
assign CPM[7155] = 12'b111111111111;
assign CPM[7156] = 12'b111111111111;
assign CPM[7157] = 12'b111111111111;
assign CPM[7158] = 12'b111111111111;
assign CPM[7159] = 12'b111111111111;
assign CPM[7160] = 12'b111111111111;
assign CPM[7161] = 12'b111111111111;
assign CPM[7162] = 12'b111111111111;
assign CPM[7163] = 12'b111111111111;
assign CPM[7164] = 12'b111111111111;
assign CPM[7165] = 12'b111111111111;
assign CPM[7166] = 12'b111111111111;
assign CPM[7167] = 12'b111111111111;
assign CPM[7168] = 12'b111111111111;
assign CPM[7169] = 12'b111111111111;
assign CPM[7170] = 12'b111111111111;
assign CPM[7171] = 12'b111111111111;
assign CPM[7172] = 12'b111111111111;
assign CPM[7173] = 12'b111111111111;
assign CPM[7174] = 12'b111111111111;
assign CPM[7175] = 12'b111111111111;
assign CPM[7176] = 12'b111111111111;
assign CPM[7177] = 12'b111111111111;
assign CPM[7178] = 12'b111111111111;
assign CPM[7179] = 12'b111111111111;
assign CPM[7180] = 12'b111111111111;
assign CPM[7181] = 12'b111111111111;
assign CPM[7182] = 12'b111111111111;
assign CPM[7183] = 12'b111111111111;
assign CPM[7184] = 12'b111111111111;
assign CPM[7185] = 12'b111111111111;
assign CPM[7186] = 12'b111111111111;
assign CPM[7187] = 12'b111111111111;
assign CPM[7188] = 12'b111111111111;
assign CPM[7189] = 12'b111111111111;
assign CPM[7190] = 12'b111111111111;
assign CPM[7191] = 12'b111111111111;
assign CPM[7192] = 12'b111111111111;
assign CPM[7193] = 12'b111111111111;
assign CPM[7194] = 12'b111111111111;
assign CPM[7195] = 12'b111111111111;
assign CPM[7196] = 12'b111111111111;
assign CPM[7197] = 12'b111111111111;
assign CPM[7198] = 12'b111111111111;
assign CPM[7199] = 12'b111111111111;
assign CPM[7200] = 12'b111111111111;
assign CPM[7201] = 12'b111111111111;
assign CPM[7202] = 12'b111111111111;
assign CPM[7203] = 12'b111111111111;
assign CPM[7204] = 12'b111111111111;
assign CPM[7205] = 12'b111111111111;
assign CPM[7206] = 12'b111111111111;
assign CPM[7207] = 12'b111111111111;
assign CPM[7208] = 12'b111111111111;
assign CPM[7209] = 12'b111111111111;
assign CPM[7210] = 12'b111111111111;
assign CPM[7211] = 12'b111111111111;
assign CPM[7212] = 12'b111111111111;
assign CPM[7213] = 12'b111111111111;
assign CPM[7214] = 12'b111111111111;
assign CPM[7215] = 12'b111111111111;
assign CPM[7216] = 12'b111111111111;
assign CPM[7217] = 12'b111111111111;
assign CPM[7218] = 12'b111111111111;
assign CPM[7219] = 12'b111111111111;
assign CPM[7220] = 12'b111111111111;
assign CPM[7221] = 12'b111111111111;
assign CPM[7222] = 12'b111111111111;
assign CPM[7223] = 12'b111111111111;
assign CPM[7224] = 12'b111111111111;
assign CPM[7225] = 12'b111111111111;
assign CPM[7226] = 12'b111111111111;
assign CPM[7227] = 12'b111111111111;
assign CPM[7228] = 12'b111111111111;
assign CPM[7229] = 12'b111111111111;
assign CPM[7230] = 12'b111111111111;
assign CPM[7231] = 12'b111111111111;
assign CPM[7232] = 12'b111111111111;
assign CPM[7233] = 12'b111111111111;
assign CPM[7234] = 12'b111111111111;
assign CPM[7235] = 12'b111111111111;
assign CPM[7236] = 12'b111111111111;
assign CPM[7237] = 12'b111111111111;
assign CPM[7238] = 12'b111111111111;
assign CPM[7239] = 12'b111111111111;
assign CPM[7240] = 12'b111111111111;
assign CPM[7241] = 12'b111111111111;
assign CPM[7242] = 12'b111111111111;
assign CPM[7243] = 12'b111111111111;
assign CPM[7244] = 12'b111111111111;
assign CPM[7245] = 12'b111111111111;
assign CPM[7246] = 12'b111111111111;
assign CPM[7247] = 12'b111111111111;
assign CPM[7248] = 12'b111111111111;
assign CPM[7249] = 12'b000000000000;
assign CPM[7250] = 12'b000000000000;
assign CPM[7251] = 12'b000000000000;
assign CPM[7252] = 12'b000000000000;
assign CPM[7253] = 12'b111111111111;
assign CPM[7254] = 12'b111111111111;
assign CPM[7255] = 12'b111111111111;
assign CPM[7256] = 12'b111111111111;
assign CPM[7257] = 12'b111111111111;
assign CPM[7258] = 12'b111111111111;
assign CPM[7259] = 12'b111111111111;
assign CPM[7260] = 12'b111111111111;
assign CPM[7261] = 12'b111111111111;
assign CPM[7262] = 12'b111111111111;
assign CPM[7263] = 12'b111111111111;
assign CPM[7264] = 12'b111111111111;
assign CPM[7265] = 12'b111111111111;
assign CPM[7266] = 12'b111111111111;
assign CPM[7267] = 12'b111111111111;
assign CPM[7268] = 12'b111111111111;
assign CPM[7269] = 12'b111111111111;
assign CPM[7270] = 12'b111111111111;
assign CPM[7271] = 12'b111111111111;
assign CPM[7272] = 12'b111111111111;
assign CPM[7273] = 12'b111111111111;
assign CPM[7274] = 12'b111111111111;
assign CPM[7275] = 12'b111111111111;
assign CPM[7276] = 12'b111111111111;
assign CPM[7277] = 12'b111111111111;
assign CPM[7278] = 12'b111111111111;
assign CPM[7279] = 12'b111111111111;
assign CPM[7280] = 12'b111111111111;
assign CPM[7281] = 12'b000000000000;
assign CPM[7282] = 12'b000000000000;
assign CPM[7283] = 12'b000000000000;
assign CPM[7284] = 12'b000000000000;
assign CPM[7285] = 12'b111111111111;
assign CPM[7286] = 12'b111111111111;
assign CPM[7287] = 12'b111111111111;
assign CPM[7288] = 12'b111111111111;
assign CPM[7289] = 12'b111111111111;
assign CPM[7290] = 12'b111111111111;
assign CPM[7291] = 12'b111111111111;
assign CPM[7292] = 12'b111111111111;
assign CPM[7293] = 12'b111111111111;
assign CPM[7294] = 12'b111111111111;
assign CPM[7295] = 12'b111111111111;
assign CPM[7296] = 12'b111111111111;
assign CPM[7297] = 12'b111111111111;
assign CPM[7298] = 12'b111111111111;
assign CPM[7299] = 12'b111111111111;
assign CPM[7300] = 12'b111111111111;
assign CPM[7301] = 12'b111111111111;
assign CPM[7302] = 12'b111111111111;
assign CPM[7303] = 12'b111111111111;
assign CPM[7304] = 12'b111111111111;
assign CPM[7305] = 12'b111111111111;
assign CPM[7306] = 12'b111111111111;
assign CPM[7307] = 12'b111111111111;
assign CPM[7308] = 12'b111111111111;
assign CPM[7309] = 12'b111111111111;
assign CPM[7310] = 12'b000000000000;
assign CPM[7311] = 12'b000000000000;
assign CPM[7312] = 12'b000000000000;
assign CPM[7313] = 12'b000000000000;
assign CPM[7314] = 12'b000000000000;
assign CPM[7315] = 12'b000000000000;
assign CPM[7316] = 12'b000000000000;
assign CPM[7317] = 12'b111111111111;
assign CPM[7318] = 12'b111111111111;
assign CPM[7319] = 12'b111111111111;
assign CPM[7320] = 12'b111111111111;
assign CPM[7321] = 12'b111111111111;
assign CPM[7322] = 12'b111111111111;
assign CPM[7323] = 12'b111111111111;
assign CPM[7324] = 12'b111111111111;
assign CPM[7325] = 12'b111111111111;
assign CPM[7326] = 12'b111111111111;
assign CPM[7327] = 12'b111111111111;
assign CPM[7328] = 12'b111111111111;
assign CPM[7329] = 12'b111111111111;
assign CPM[7330] = 12'b111111111111;
assign CPM[7331] = 12'b111111111111;
assign CPM[7332] = 12'b111111111111;
assign CPM[7333] = 12'b111111111111;
assign CPM[7334] = 12'b111111111111;
assign CPM[7335] = 12'b111111111111;
assign CPM[7336] = 12'b111111111111;
assign CPM[7337] = 12'b111111111111;
assign CPM[7338] = 12'b111111111111;
assign CPM[7339] = 12'b111111111111;
assign CPM[7340] = 12'b111111111111;
assign CPM[7341] = 12'b111111111111;
assign CPM[7342] = 12'b000000000000;
assign CPM[7343] = 12'b000000000000;
assign CPM[7344] = 12'b000000000000;
assign CPM[7345] = 12'b000000000000;
assign CPM[7346] = 12'b000000000000;
assign CPM[7347] = 12'b000000000000;
assign CPM[7348] = 12'b000000000000;
assign CPM[7349] = 12'b111111111111;
assign CPM[7350] = 12'b111111111111;
assign CPM[7351] = 12'b111111111111;
assign CPM[7352] = 12'b111111111111;
assign CPM[7353] = 12'b111111111111;
assign CPM[7354] = 12'b111111111111;
assign CPM[7355] = 12'b111111111111;
assign CPM[7356] = 12'b111111111111;
assign CPM[7357] = 12'b111111111111;
assign CPM[7358] = 12'b111111111111;
assign CPM[7359] = 12'b111111111111;
assign CPM[7360] = 12'b111111111111;
assign CPM[7361] = 12'b111111111111;
assign CPM[7362] = 12'b111111111111;
assign CPM[7363] = 12'b111111111111;
assign CPM[7364] = 12'b111111111111;
assign CPM[7365] = 12'b111111111111;
assign CPM[7366] = 12'b111111111111;
assign CPM[7367] = 12'b111111111111;
assign CPM[7368] = 12'b111111111111;
assign CPM[7369] = 12'b111111111111;
assign CPM[7370] = 12'b111111111111;
assign CPM[7371] = 12'b111111111111;
assign CPM[7372] = 12'b111111111111;
assign CPM[7373] = 12'b111111111111;
assign CPM[7374] = 12'b000000000000;
assign CPM[7375] = 12'b000000000000;
assign CPM[7376] = 12'b000000000000;
assign CPM[7377] = 12'b000000000000;
assign CPM[7378] = 12'b000000000000;
assign CPM[7379] = 12'b000000000000;
assign CPM[7380] = 12'b000000000000;
assign CPM[7381] = 12'b111111111111;
assign CPM[7382] = 12'b111111111111;
assign CPM[7383] = 12'b111111111111;
assign CPM[7384] = 12'b111111111111;
assign CPM[7385] = 12'b111111111111;
assign CPM[7386] = 12'b111111111111;
assign CPM[7387] = 12'b111111111111;
assign CPM[7388] = 12'b111111111111;
assign CPM[7389] = 12'b111111111111;
assign CPM[7390] = 12'b111111111111;
assign CPM[7391] = 12'b111111111111;
assign CPM[7392] = 12'b111111111111;
assign CPM[7393] = 12'b111111111111;
assign CPM[7394] = 12'b111111111111;
assign CPM[7395] = 12'b111111111111;
assign CPM[7396] = 12'b111111111111;
assign CPM[7397] = 12'b111111111111;
assign CPM[7398] = 12'b111111111111;
assign CPM[7399] = 12'b111111111111;
assign CPM[7400] = 12'b111111111111;
assign CPM[7401] = 12'b111111111111;
assign CPM[7402] = 12'b111111111111;
assign CPM[7403] = 12'b111111111111;
assign CPM[7404] = 12'b111111111111;
assign CPM[7405] = 12'b111111111111;
assign CPM[7406] = 12'b000000000000;
assign CPM[7407] = 12'b000000000000;
assign CPM[7408] = 12'b000000000000;
assign CPM[7409] = 12'b000000000000;
assign CPM[7410] = 12'b000000000000;
assign CPM[7411] = 12'b000000000000;
assign CPM[7412] = 12'b000000000000;
assign CPM[7413] = 12'b111111111111;
assign CPM[7414] = 12'b111111111111;
assign CPM[7415] = 12'b111111111111;
assign CPM[7416] = 12'b111111111111;
assign CPM[7417] = 12'b111111111111;
assign CPM[7418] = 12'b111111111111;
assign CPM[7419] = 12'b111111111111;
assign CPM[7420] = 12'b111111111111;
assign CPM[7421] = 12'b111111111111;
assign CPM[7422] = 12'b111111111111;
assign CPM[7423] = 12'b111111111111;
assign CPM[7424] = 12'b111111111111;
assign CPM[7425] = 12'b111111111111;
assign CPM[7426] = 12'b111111111111;
assign CPM[7427] = 12'b111111111111;
assign CPM[7428] = 12'b111111111111;
assign CPM[7429] = 12'b111111111111;
assign CPM[7430] = 12'b111111111111;
assign CPM[7431] = 12'b111111111111;
assign CPM[7432] = 12'b111111111111;
assign CPM[7433] = 12'b111111111111;
assign CPM[7434] = 12'b111111111111;
assign CPM[7435] = 12'b000000000000;
assign CPM[7436] = 12'b000000000000;
assign CPM[7437] = 12'b000000000000;
assign CPM[7438] = 12'b000000000000;
assign CPM[7439] = 12'b111111111111;
assign CPM[7440] = 12'b111111111111;
assign CPM[7441] = 12'b000000000000;
assign CPM[7442] = 12'b000000000000;
assign CPM[7443] = 12'b000000000000;
assign CPM[7444] = 12'b000000000000;
assign CPM[7445] = 12'b111111111111;
assign CPM[7446] = 12'b111111111111;
assign CPM[7447] = 12'b111111111111;
assign CPM[7448] = 12'b111111111111;
assign CPM[7449] = 12'b111111111111;
assign CPM[7450] = 12'b111111111111;
assign CPM[7451] = 12'b111111111111;
assign CPM[7452] = 12'b111111111111;
assign CPM[7453] = 12'b111111111111;
assign CPM[7454] = 12'b111111111111;
assign CPM[7455] = 12'b111111111111;
assign CPM[7456] = 12'b111111111111;
assign CPM[7457] = 12'b111111111111;
assign CPM[7458] = 12'b111111111111;
assign CPM[7459] = 12'b111111111111;
assign CPM[7460] = 12'b111111111111;
assign CPM[7461] = 12'b111111111111;
assign CPM[7462] = 12'b111111111111;
assign CPM[7463] = 12'b111111111111;
assign CPM[7464] = 12'b111111111111;
assign CPM[7465] = 12'b111111111111;
assign CPM[7466] = 12'b111111111111;
assign CPM[7467] = 12'b000000000000;
assign CPM[7468] = 12'b000000000000;
assign CPM[7469] = 12'b000000000000;
assign CPM[7470] = 12'b000000000000;
assign CPM[7471] = 12'b111111111111;
assign CPM[7472] = 12'b111111111111;
assign CPM[7473] = 12'b000000000000;
assign CPM[7474] = 12'b000000000000;
assign CPM[7475] = 12'b000000000000;
assign CPM[7476] = 12'b000000000000;
assign CPM[7477] = 12'b111111111111;
assign CPM[7478] = 12'b111111111111;
assign CPM[7479] = 12'b111111111111;
assign CPM[7480] = 12'b111111111111;
assign CPM[7481] = 12'b111111111111;
assign CPM[7482] = 12'b111111111111;
assign CPM[7483] = 12'b111111111111;
assign CPM[7484] = 12'b111111111111;
assign CPM[7485] = 12'b111111111111;
assign CPM[7486] = 12'b111111111111;
assign CPM[7487] = 12'b111111111111;
assign CPM[7488] = 12'b111111111111;
assign CPM[7489] = 12'b111111111111;
assign CPM[7490] = 12'b111111111111;
assign CPM[7491] = 12'b111111111111;
assign CPM[7492] = 12'b111111111111;
assign CPM[7493] = 12'b111111111111;
assign CPM[7494] = 12'b111111111111;
assign CPM[7495] = 12'b111111111111;
assign CPM[7496] = 12'b111111111111;
assign CPM[7497] = 12'b111111111111;
assign CPM[7498] = 12'b111111111111;
assign CPM[7499] = 12'b000000000000;
assign CPM[7500] = 12'b000000000000;
assign CPM[7501] = 12'b000000000000;
assign CPM[7502] = 12'b000000000000;
assign CPM[7503] = 12'b111111111111;
assign CPM[7504] = 12'b111111111111;
assign CPM[7505] = 12'b000000000000;
assign CPM[7506] = 12'b000000000000;
assign CPM[7507] = 12'b000000000000;
assign CPM[7508] = 12'b000000000000;
assign CPM[7509] = 12'b111111111111;
assign CPM[7510] = 12'b111111111111;
assign CPM[7511] = 12'b111111111111;
assign CPM[7512] = 12'b111111111111;
assign CPM[7513] = 12'b111111111111;
assign CPM[7514] = 12'b111111111111;
assign CPM[7515] = 12'b111111111111;
assign CPM[7516] = 12'b111111111111;
assign CPM[7517] = 12'b111111111111;
assign CPM[7518] = 12'b111111111111;
assign CPM[7519] = 12'b111111111111;
assign CPM[7520] = 12'b111111111111;
assign CPM[7521] = 12'b111111111111;
assign CPM[7522] = 12'b111111111111;
assign CPM[7523] = 12'b111111111111;
assign CPM[7524] = 12'b111111111111;
assign CPM[7525] = 12'b111111111111;
assign CPM[7526] = 12'b111111111111;
assign CPM[7527] = 12'b111111111111;
assign CPM[7528] = 12'b111111111111;
assign CPM[7529] = 12'b111111111111;
assign CPM[7530] = 12'b111111111111;
assign CPM[7531] = 12'b000000000000;
assign CPM[7532] = 12'b000000000000;
assign CPM[7533] = 12'b000000000000;
assign CPM[7534] = 12'b000000000000;
assign CPM[7535] = 12'b111111111111;
assign CPM[7536] = 12'b111111111111;
assign CPM[7537] = 12'b000000000000;
assign CPM[7538] = 12'b000000000000;
assign CPM[7539] = 12'b000000000000;
assign CPM[7540] = 12'b000000000000;
assign CPM[7541] = 12'b111111111111;
assign CPM[7542] = 12'b111111111111;
assign CPM[7543] = 12'b111111111111;
assign CPM[7544] = 12'b111111111111;
assign CPM[7545] = 12'b111111111111;
assign CPM[7546] = 12'b111111111111;
assign CPM[7547] = 12'b111111111111;
assign CPM[7548] = 12'b111111111111;
assign CPM[7549] = 12'b111111111111;
assign CPM[7550] = 12'b111111111111;
assign CPM[7551] = 12'b111111111111;
assign CPM[7552] = 12'b111111111111;
assign CPM[7553] = 12'b111111111111;
assign CPM[7554] = 12'b111111111111;
assign CPM[7555] = 12'b111111111111;
assign CPM[7556] = 12'b111111111111;
assign CPM[7557] = 12'b111111111111;
assign CPM[7558] = 12'b111111111111;
assign CPM[7559] = 12'b111111111111;
assign CPM[7560] = 12'b000000000000;
assign CPM[7561] = 12'b000000000000;
assign CPM[7562] = 12'b000000000000;
assign CPM[7563] = 12'b000000000000;
assign CPM[7564] = 12'b111111111111;
assign CPM[7565] = 12'b111111111111;
assign CPM[7566] = 12'b111111111111;
assign CPM[7567] = 12'b111111111111;
assign CPM[7568] = 12'b111111111111;
assign CPM[7569] = 12'b000000000000;
assign CPM[7570] = 12'b000000000000;
assign CPM[7571] = 12'b000000000000;
assign CPM[7572] = 12'b000000000000;
assign CPM[7573] = 12'b111111111111;
assign CPM[7574] = 12'b111111111111;
assign CPM[7575] = 12'b111111111111;
assign CPM[7576] = 12'b111111111111;
assign CPM[7577] = 12'b111111111111;
assign CPM[7578] = 12'b111111111111;
assign CPM[7579] = 12'b111111111111;
assign CPM[7580] = 12'b111111111111;
assign CPM[7581] = 12'b111111111111;
assign CPM[7582] = 12'b111111111111;
assign CPM[7583] = 12'b111111111111;
assign CPM[7584] = 12'b111111111111;
assign CPM[7585] = 12'b111111111111;
assign CPM[7586] = 12'b111111111111;
assign CPM[7587] = 12'b111111111111;
assign CPM[7588] = 12'b111111111111;
assign CPM[7589] = 12'b111111111111;
assign CPM[7590] = 12'b111111111111;
assign CPM[7591] = 12'b111111111111;
assign CPM[7592] = 12'b000000000000;
assign CPM[7593] = 12'b000000000000;
assign CPM[7594] = 12'b000000000000;
assign CPM[7595] = 12'b000000000000;
assign CPM[7596] = 12'b111111111111;
assign CPM[7597] = 12'b111111111111;
assign CPM[7598] = 12'b111111111111;
assign CPM[7599] = 12'b111111111111;
assign CPM[7600] = 12'b111111111111;
assign CPM[7601] = 12'b000000000000;
assign CPM[7602] = 12'b000000000000;
assign CPM[7603] = 12'b000000000000;
assign CPM[7604] = 12'b000000000000;
assign CPM[7605] = 12'b111111111111;
assign CPM[7606] = 12'b111111111111;
assign CPM[7607] = 12'b111111111111;
assign CPM[7608] = 12'b111111111111;
assign CPM[7609] = 12'b111111111111;
assign CPM[7610] = 12'b111111111111;
assign CPM[7611] = 12'b111111111111;
assign CPM[7612] = 12'b111111111111;
assign CPM[7613] = 12'b111111111111;
assign CPM[7614] = 12'b111111111111;
assign CPM[7615] = 12'b111111111111;
assign CPM[7616] = 12'b111111111111;
assign CPM[7617] = 12'b111111111111;
assign CPM[7618] = 12'b111111111111;
assign CPM[7619] = 12'b111111111111;
assign CPM[7620] = 12'b111111111111;
assign CPM[7621] = 12'b111111111111;
assign CPM[7622] = 12'b111111111111;
assign CPM[7623] = 12'b111111111111;
assign CPM[7624] = 12'b000000000000;
assign CPM[7625] = 12'b000000000000;
assign CPM[7626] = 12'b000000000000;
assign CPM[7627] = 12'b000000000000;
assign CPM[7628] = 12'b111111111111;
assign CPM[7629] = 12'b111111111111;
assign CPM[7630] = 12'b111111111111;
assign CPM[7631] = 12'b111111111111;
assign CPM[7632] = 12'b111111111111;
assign CPM[7633] = 12'b000000000000;
assign CPM[7634] = 12'b000000000000;
assign CPM[7635] = 12'b000000000000;
assign CPM[7636] = 12'b000000000000;
assign CPM[7637] = 12'b111111111111;
assign CPM[7638] = 12'b111111111111;
assign CPM[7639] = 12'b111111111111;
assign CPM[7640] = 12'b111111111111;
assign CPM[7641] = 12'b111111111111;
assign CPM[7642] = 12'b111111111111;
assign CPM[7643] = 12'b111111111111;
assign CPM[7644] = 12'b111111111111;
assign CPM[7645] = 12'b111111111111;
assign CPM[7646] = 12'b111111111111;
assign CPM[7647] = 12'b111111111111;
assign CPM[7648] = 12'b111111111111;
assign CPM[7649] = 12'b111111111111;
assign CPM[7650] = 12'b111111111111;
assign CPM[7651] = 12'b111111111111;
assign CPM[7652] = 12'b111111111111;
assign CPM[7653] = 12'b111111111111;
assign CPM[7654] = 12'b111111111111;
assign CPM[7655] = 12'b111111111111;
assign CPM[7656] = 12'b000000000000;
assign CPM[7657] = 12'b000000000000;
assign CPM[7658] = 12'b000000000000;
assign CPM[7659] = 12'b000000000000;
assign CPM[7660] = 12'b111111111111;
assign CPM[7661] = 12'b111111111111;
assign CPM[7662] = 12'b111111111111;
assign CPM[7663] = 12'b111111111111;
assign CPM[7664] = 12'b111111111111;
assign CPM[7665] = 12'b000000000000;
assign CPM[7666] = 12'b000000000000;
assign CPM[7667] = 12'b000000000000;
assign CPM[7668] = 12'b000000000000;
assign CPM[7669] = 12'b111111111111;
assign CPM[7670] = 12'b111111111111;
assign CPM[7671] = 12'b111111111111;
assign CPM[7672] = 12'b111111111111;
assign CPM[7673] = 12'b111111111111;
assign CPM[7674] = 12'b111111111111;
assign CPM[7675] = 12'b111111111111;
assign CPM[7676] = 12'b111111111111;
assign CPM[7677] = 12'b111111111111;
assign CPM[7678] = 12'b111111111111;
assign CPM[7679] = 12'b111111111111;
assign CPM[7680] = 12'b111111111111;
assign CPM[7681] = 12'b111111111111;
assign CPM[7682] = 12'b111111111111;
assign CPM[7683] = 12'b111111111111;
assign CPM[7684] = 12'b111111111111;
assign CPM[7685] = 12'b000000000000;
assign CPM[7686] = 12'b000000000000;
assign CPM[7687] = 12'b000000000000;
assign CPM[7688] = 12'b000000000000;
assign CPM[7689] = 12'b111111111111;
assign CPM[7690] = 12'b111111111111;
assign CPM[7691] = 12'b111111111111;
assign CPM[7692] = 12'b111111111111;
assign CPM[7693] = 12'b111111111111;
assign CPM[7694] = 12'b111111111111;
assign CPM[7695] = 12'b111111111111;
assign CPM[7696] = 12'b111111111111;
assign CPM[7697] = 12'b000000000000;
assign CPM[7698] = 12'b000000000000;
assign CPM[7699] = 12'b000000000000;
assign CPM[7700] = 12'b000000000000;
assign CPM[7701] = 12'b111111111111;
assign CPM[7702] = 12'b111111111111;
assign CPM[7703] = 12'b111111111111;
assign CPM[7704] = 12'b111111111111;
assign CPM[7705] = 12'b111111111111;
assign CPM[7706] = 12'b111111111111;
assign CPM[7707] = 12'b111111111111;
assign CPM[7708] = 12'b111111111111;
assign CPM[7709] = 12'b111111111111;
assign CPM[7710] = 12'b111111111111;
assign CPM[7711] = 12'b111111111111;
assign CPM[7712] = 12'b111111111111;
assign CPM[7713] = 12'b111111111111;
assign CPM[7714] = 12'b111111111111;
assign CPM[7715] = 12'b111111111111;
assign CPM[7716] = 12'b111111111111;
assign CPM[7717] = 12'b000000000000;
assign CPM[7718] = 12'b000000000000;
assign CPM[7719] = 12'b000000000000;
assign CPM[7720] = 12'b000000000000;
assign CPM[7721] = 12'b111111111111;
assign CPM[7722] = 12'b111111111111;
assign CPM[7723] = 12'b111111111111;
assign CPM[7724] = 12'b111111111111;
assign CPM[7725] = 12'b111111111111;
assign CPM[7726] = 12'b111111111111;
assign CPM[7727] = 12'b111111111111;
assign CPM[7728] = 12'b111111111111;
assign CPM[7729] = 12'b000000000000;
assign CPM[7730] = 12'b000000000000;
assign CPM[7731] = 12'b000000000000;
assign CPM[7732] = 12'b000000000000;
assign CPM[7733] = 12'b111111111111;
assign CPM[7734] = 12'b111111111111;
assign CPM[7735] = 12'b111111111111;
assign CPM[7736] = 12'b111111111111;
assign CPM[7737] = 12'b111111111111;
assign CPM[7738] = 12'b111111111111;
assign CPM[7739] = 12'b111111111111;
assign CPM[7740] = 12'b111111111111;
assign CPM[7741] = 12'b111111111111;
assign CPM[7742] = 12'b111111111111;
assign CPM[7743] = 12'b111111111111;
assign CPM[7744] = 12'b111111111111;
assign CPM[7745] = 12'b111111111111;
assign CPM[7746] = 12'b111111111111;
assign CPM[7747] = 12'b111111111111;
assign CPM[7748] = 12'b111111111111;
assign CPM[7749] = 12'b000000000000;
assign CPM[7750] = 12'b000000000000;
assign CPM[7751] = 12'b000000000000;
assign CPM[7752] = 12'b000000000000;
assign CPM[7753] = 12'b111111111111;
assign CPM[7754] = 12'b111111111111;
assign CPM[7755] = 12'b111111111111;
assign CPM[7756] = 12'b111111111111;
assign CPM[7757] = 12'b111111111111;
assign CPM[7758] = 12'b111111111111;
assign CPM[7759] = 12'b111111111111;
assign CPM[7760] = 12'b111111111111;
assign CPM[7761] = 12'b000000000000;
assign CPM[7762] = 12'b000000000000;
assign CPM[7763] = 12'b000000000000;
assign CPM[7764] = 12'b000000000000;
assign CPM[7765] = 12'b111111111111;
assign CPM[7766] = 12'b111111111111;
assign CPM[7767] = 12'b111111111111;
assign CPM[7768] = 12'b111111111111;
assign CPM[7769] = 12'b111111111111;
assign CPM[7770] = 12'b111111111111;
assign CPM[7771] = 12'b111111111111;
assign CPM[7772] = 12'b111111111111;
assign CPM[7773] = 12'b111111111111;
assign CPM[7774] = 12'b111111111111;
assign CPM[7775] = 12'b111111111111;
assign CPM[7776] = 12'b111111111111;
assign CPM[7777] = 12'b111111111111;
assign CPM[7778] = 12'b111111111111;
assign CPM[7779] = 12'b111111111111;
assign CPM[7780] = 12'b111111111111;
assign CPM[7781] = 12'b000000000000;
assign CPM[7782] = 12'b000000000000;
assign CPM[7783] = 12'b000000000000;
assign CPM[7784] = 12'b000000000000;
assign CPM[7785] = 12'b000000000000;
assign CPM[7786] = 12'b000000000000;
assign CPM[7787] = 12'b000000000000;
assign CPM[7788] = 12'b000000000000;
assign CPM[7789] = 12'b000000000000;
assign CPM[7790] = 12'b000000000000;
assign CPM[7791] = 12'b000000000000;
assign CPM[7792] = 12'b000000000000;
assign CPM[7793] = 12'b000000000000;
assign CPM[7794] = 12'b000000000000;
assign CPM[7795] = 12'b000000000000;
assign CPM[7796] = 12'b000000000000;
assign CPM[7797] = 12'b000000000000;
assign CPM[7798] = 12'b000000000000;
assign CPM[7799] = 12'b000000000000;
assign CPM[7800] = 12'b000000000000;
assign CPM[7801] = 12'b000000000000;
assign CPM[7802] = 12'b111111111111;
assign CPM[7803] = 12'b111111111111;
assign CPM[7804] = 12'b111111111111;
assign CPM[7805] = 12'b111111111111;
assign CPM[7806] = 12'b111111111111;
assign CPM[7807] = 12'b111111111111;
assign CPM[7808] = 12'b111111111111;
assign CPM[7809] = 12'b111111111111;
assign CPM[7810] = 12'b111111111111;
assign CPM[7811] = 12'b111111111111;
assign CPM[7812] = 12'b111111111111;
assign CPM[7813] = 12'b000000000000;
assign CPM[7814] = 12'b000000000000;
assign CPM[7815] = 12'b000000000000;
assign CPM[7816] = 12'b000000000000;
assign CPM[7817] = 12'b000000000000;
assign CPM[7818] = 12'b000000000000;
assign CPM[7819] = 12'b000000000000;
assign CPM[7820] = 12'b000000000000;
assign CPM[7821] = 12'b000000000000;
assign CPM[7822] = 12'b000000000000;
assign CPM[7823] = 12'b000000000000;
assign CPM[7824] = 12'b000000000000;
assign CPM[7825] = 12'b000000000000;
assign CPM[7826] = 12'b000000000000;
assign CPM[7827] = 12'b000000000000;
assign CPM[7828] = 12'b000000000000;
assign CPM[7829] = 12'b000000000000;
assign CPM[7830] = 12'b000000000000;
assign CPM[7831] = 12'b000000000000;
assign CPM[7832] = 12'b000000000000;
assign CPM[7833] = 12'b000000000000;
assign CPM[7834] = 12'b111111111111;
assign CPM[7835] = 12'b111111111111;
assign CPM[7836] = 12'b111111111111;
assign CPM[7837] = 12'b111111111111;
assign CPM[7838] = 12'b111111111111;
assign CPM[7839] = 12'b111111111111;
assign CPM[7840] = 12'b111111111111;
assign CPM[7841] = 12'b111111111111;
assign CPM[7842] = 12'b111111111111;
assign CPM[7843] = 12'b111111111111;
assign CPM[7844] = 12'b111111111111;
assign CPM[7845] = 12'b000000000000;
assign CPM[7846] = 12'b000000000000;
assign CPM[7847] = 12'b000000000000;
assign CPM[7848] = 12'b000000000000;
assign CPM[7849] = 12'b000000000000;
assign CPM[7850] = 12'b000000000000;
assign CPM[7851] = 12'b000000000000;
assign CPM[7852] = 12'b000000000000;
assign CPM[7853] = 12'b000000000000;
assign CPM[7854] = 12'b000000000000;
assign CPM[7855] = 12'b000000000000;
assign CPM[7856] = 12'b000000000000;
assign CPM[7857] = 12'b000000000000;
assign CPM[7858] = 12'b000000000000;
assign CPM[7859] = 12'b000000000000;
assign CPM[7860] = 12'b000000000000;
assign CPM[7861] = 12'b000000000000;
assign CPM[7862] = 12'b000000000000;
assign CPM[7863] = 12'b000000000000;
assign CPM[7864] = 12'b000000000000;
assign CPM[7865] = 12'b000000000000;
assign CPM[7866] = 12'b111111111111;
assign CPM[7867] = 12'b111111111111;
assign CPM[7868] = 12'b111111111111;
assign CPM[7869] = 12'b111111111111;
assign CPM[7870] = 12'b111111111111;
assign CPM[7871] = 12'b111111111111;
assign CPM[7872] = 12'b111111111111;
assign CPM[7873] = 12'b111111111111;
assign CPM[7874] = 12'b111111111111;
assign CPM[7875] = 12'b111111111111;
assign CPM[7876] = 12'b111111111111;
assign CPM[7877] = 12'b000000000000;
assign CPM[7878] = 12'b000000000000;
assign CPM[7879] = 12'b000000000000;
assign CPM[7880] = 12'b000000000000;
assign CPM[7881] = 12'b000000000000;
assign CPM[7882] = 12'b000000000000;
assign CPM[7883] = 12'b000000000000;
assign CPM[7884] = 12'b000000000000;
assign CPM[7885] = 12'b000000000000;
assign CPM[7886] = 12'b000000000000;
assign CPM[7887] = 12'b000000000000;
assign CPM[7888] = 12'b000000000000;
assign CPM[7889] = 12'b000000000000;
assign CPM[7890] = 12'b000000000000;
assign CPM[7891] = 12'b000000000000;
assign CPM[7892] = 12'b000000000000;
assign CPM[7893] = 12'b000000000000;
assign CPM[7894] = 12'b000000000000;
assign CPM[7895] = 12'b000000000000;
assign CPM[7896] = 12'b000000000000;
assign CPM[7897] = 12'b000000000000;
assign CPM[7898] = 12'b111111111111;
assign CPM[7899] = 12'b111111111111;
assign CPM[7900] = 12'b111111111111;
assign CPM[7901] = 12'b111111111111;
assign CPM[7902] = 12'b111111111111;
assign CPM[7903] = 12'b111111111111;
assign CPM[7904] = 12'b111111111111;
assign CPM[7905] = 12'b111111111111;
assign CPM[7906] = 12'b111111111111;
assign CPM[7907] = 12'b111111111111;
assign CPM[7908] = 12'b111111111111;
assign CPM[7909] = 12'b111111111111;
assign CPM[7910] = 12'b111111111111;
assign CPM[7911] = 12'b111111111111;
assign CPM[7912] = 12'b111111111111;
assign CPM[7913] = 12'b111111111111;
assign CPM[7914] = 12'b111111111111;
assign CPM[7915] = 12'b111111111111;
assign CPM[7916] = 12'b111111111111;
assign CPM[7917] = 12'b111111111111;
assign CPM[7918] = 12'b111111111111;
assign CPM[7919] = 12'b111111111111;
assign CPM[7920] = 12'b111111111111;
assign CPM[7921] = 12'b000000000000;
assign CPM[7922] = 12'b000000000000;
assign CPM[7923] = 12'b000000000000;
assign CPM[7924] = 12'b000000000000;
assign CPM[7925] = 12'b111111111111;
assign CPM[7926] = 12'b111111111111;
assign CPM[7927] = 12'b111111111111;
assign CPM[7928] = 12'b111111111111;
assign CPM[7929] = 12'b111111111111;
assign CPM[7930] = 12'b111111111111;
assign CPM[7931] = 12'b111111111111;
assign CPM[7932] = 12'b111111111111;
assign CPM[7933] = 12'b111111111111;
assign CPM[7934] = 12'b111111111111;
assign CPM[7935] = 12'b111111111111;
assign CPM[7936] = 12'b111111111111;
assign CPM[7937] = 12'b111111111111;
assign CPM[7938] = 12'b111111111111;
assign CPM[7939] = 12'b111111111111;
assign CPM[7940] = 12'b111111111111;
assign CPM[7941] = 12'b111111111111;
assign CPM[7942] = 12'b111111111111;
assign CPM[7943] = 12'b111111111111;
assign CPM[7944] = 12'b111111111111;
assign CPM[7945] = 12'b111111111111;
assign CPM[7946] = 12'b111111111111;
assign CPM[7947] = 12'b111111111111;
assign CPM[7948] = 12'b111111111111;
assign CPM[7949] = 12'b111111111111;
assign CPM[7950] = 12'b111111111111;
assign CPM[7951] = 12'b111111111111;
assign CPM[7952] = 12'b111111111111;
assign CPM[7953] = 12'b000000000000;
assign CPM[7954] = 12'b000000000000;
assign CPM[7955] = 12'b000000000000;
assign CPM[7956] = 12'b000000000000;
assign CPM[7957] = 12'b111111111111;
assign CPM[7958] = 12'b111111111111;
assign CPM[7959] = 12'b111111111111;
assign CPM[7960] = 12'b111111111111;
assign CPM[7961] = 12'b111111111111;
assign CPM[7962] = 12'b111111111111;
assign CPM[7963] = 12'b111111111111;
assign CPM[7964] = 12'b111111111111;
assign CPM[7965] = 12'b111111111111;
assign CPM[7966] = 12'b111111111111;
assign CPM[7967] = 12'b111111111111;
assign CPM[7968] = 12'b111111111111;
assign CPM[7969] = 12'b111111111111;
assign CPM[7970] = 12'b111111111111;
assign CPM[7971] = 12'b111111111111;
assign CPM[7972] = 12'b111111111111;
assign CPM[7973] = 12'b111111111111;
assign CPM[7974] = 12'b111111111111;
assign CPM[7975] = 12'b111111111111;
assign CPM[7976] = 12'b111111111111;
assign CPM[7977] = 12'b111111111111;
assign CPM[7978] = 12'b111111111111;
assign CPM[7979] = 12'b111111111111;
assign CPM[7980] = 12'b111111111111;
assign CPM[7981] = 12'b111111111111;
assign CPM[7982] = 12'b111111111111;
assign CPM[7983] = 12'b111111111111;
assign CPM[7984] = 12'b111111111111;
assign CPM[7985] = 12'b000000000000;
assign CPM[7986] = 12'b000000000000;
assign CPM[7987] = 12'b000000000000;
assign CPM[7988] = 12'b000000000000;
assign CPM[7989] = 12'b111111111111;
assign CPM[7990] = 12'b111111111111;
assign CPM[7991] = 12'b111111111111;
assign CPM[7992] = 12'b111111111111;
assign CPM[7993] = 12'b111111111111;
assign CPM[7994] = 12'b111111111111;
assign CPM[7995] = 12'b111111111111;
assign CPM[7996] = 12'b111111111111;
assign CPM[7997] = 12'b111111111111;
assign CPM[7998] = 12'b111111111111;
assign CPM[7999] = 12'b111111111111;
assign CPM[8000] = 12'b111111111111;
assign CPM[8001] = 12'b111111111111;
assign CPM[8002] = 12'b111111111111;
assign CPM[8003] = 12'b111111111111;
assign CPM[8004] = 12'b111111111111;
assign CPM[8005] = 12'b111111111111;
assign CPM[8006] = 12'b111111111111;
assign CPM[8007] = 12'b111111111111;
assign CPM[8008] = 12'b111111111111;
assign CPM[8009] = 12'b111111111111;
assign CPM[8010] = 12'b111111111111;
assign CPM[8011] = 12'b111111111111;
assign CPM[8012] = 12'b111111111111;
assign CPM[8013] = 12'b111111111111;
assign CPM[8014] = 12'b111111111111;
assign CPM[8015] = 12'b111111111111;
assign CPM[8016] = 12'b111111111111;
assign CPM[8017] = 12'b000000000000;
assign CPM[8018] = 12'b000000000000;
assign CPM[8019] = 12'b000000000000;
assign CPM[8020] = 12'b000000000000;
assign CPM[8021] = 12'b111111111111;
assign CPM[8022] = 12'b111111111111;
assign CPM[8023] = 12'b111111111111;
assign CPM[8024] = 12'b111111111111;
assign CPM[8025] = 12'b111111111111;
assign CPM[8026] = 12'b111111111111;
assign CPM[8027] = 12'b111111111111;
assign CPM[8028] = 12'b111111111111;
assign CPM[8029] = 12'b111111111111;
assign CPM[8030] = 12'b111111111111;
assign CPM[8031] = 12'b111111111111;
assign CPM[8032] = 12'b111111111111;
assign CPM[8033] = 12'b111111111111;
assign CPM[8034] = 12'b111111111111;
assign CPM[8035] = 12'b111111111111;
assign CPM[8036] = 12'b111111111111;
assign CPM[8037] = 12'b111111111111;
assign CPM[8038] = 12'b111111111111;
assign CPM[8039] = 12'b111111111111;
assign CPM[8040] = 12'b111111111111;
assign CPM[8041] = 12'b111111111111;
assign CPM[8042] = 12'b111111111111;
assign CPM[8043] = 12'b111111111111;
assign CPM[8044] = 12'b111111111111;
assign CPM[8045] = 12'b111111111111;
assign CPM[8046] = 12'b111111111111;
assign CPM[8047] = 12'b111111111111;
assign CPM[8048] = 12'b111111111111;
assign CPM[8049] = 12'b000000000000;
assign CPM[8050] = 12'b000000000000;
assign CPM[8051] = 12'b000000000000;
assign CPM[8052] = 12'b000000000000;
assign CPM[8053] = 12'b111111111111;
assign CPM[8054] = 12'b111111111111;
assign CPM[8055] = 12'b111111111111;
assign CPM[8056] = 12'b111111111111;
assign CPM[8057] = 12'b111111111111;
assign CPM[8058] = 12'b111111111111;
assign CPM[8059] = 12'b111111111111;
assign CPM[8060] = 12'b111111111111;
assign CPM[8061] = 12'b111111111111;
assign CPM[8062] = 12'b111111111111;
assign CPM[8063] = 12'b111111111111;
assign CPM[8064] = 12'b111111111111;
assign CPM[8065] = 12'b111111111111;
assign CPM[8066] = 12'b111111111111;
assign CPM[8067] = 12'b111111111111;
assign CPM[8068] = 12'b111111111111;
assign CPM[8069] = 12'b111111111111;
assign CPM[8070] = 12'b111111111111;
assign CPM[8071] = 12'b111111111111;
assign CPM[8072] = 12'b111111111111;
assign CPM[8073] = 12'b111111111111;
assign CPM[8074] = 12'b111111111111;
assign CPM[8075] = 12'b111111111111;
assign CPM[8076] = 12'b111111111111;
assign CPM[8077] = 12'b111111111111;
assign CPM[8078] = 12'b111111111111;
assign CPM[8079] = 12'b111111111111;
assign CPM[8080] = 12'b111111111111;
assign CPM[8081] = 12'b000000000000;
assign CPM[8082] = 12'b000000000000;
assign CPM[8083] = 12'b000000000000;
assign CPM[8084] = 12'b000000000000;
assign CPM[8085] = 12'b111111111111;
assign CPM[8086] = 12'b111111111111;
assign CPM[8087] = 12'b111111111111;
assign CPM[8088] = 12'b111111111111;
assign CPM[8089] = 12'b111111111111;
assign CPM[8090] = 12'b111111111111;
assign CPM[8091] = 12'b111111111111;
assign CPM[8092] = 12'b111111111111;
assign CPM[8093] = 12'b111111111111;
assign CPM[8094] = 12'b111111111111;
assign CPM[8095] = 12'b111111111111;
assign CPM[8096] = 12'b111111111111;
assign CPM[8097] = 12'b111111111111;
assign CPM[8098] = 12'b111111111111;
assign CPM[8099] = 12'b111111111111;
assign CPM[8100] = 12'b111111111111;
assign CPM[8101] = 12'b111111111111;
assign CPM[8102] = 12'b111111111111;
assign CPM[8103] = 12'b111111111111;
assign CPM[8104] = 12'b111111111111;
assign CPM[8105] = 12'b111111111111;
assign CPM[8106] = 12'b111111111111;
assign CPM[8107] = 12'b111111111111;
assign CPM[8108] = 12'b111111111111;
assign CPM[8109] = 12'b111111111111;
assign CPM[8110] = 12'b111111111111;
assign CPM[8111] = 12'b111111111111;
assign CPM[8112] = 12'b111111111111;
assign CPM[8113] = 12'b000000000000;
assign CPM[8114] = 12'b000000000000;
assign CPM[8115] = 12'b000000000000;
assign CPM[8116] = 12'b000000000000;
assign CPM[8117] = 12'b111111111111;
assign CPM[8118] = 12'b111111111111;
assign CPM[8119] = 12'b111111111111;
assign CPM[8120] = 12'b111111111111;
assign CPM[8121] = 12'b111111111111;
assign CPM[8122] = 12'b111111111111;
assign CPM[8123] = 12'b111111111111;
assign CPM[8124] = 12'b111111111111;
assign CPM[8125] = 12'b111111111111;
assign CPM[8126] = 12'b111111111111;
assign CPM[8127] = 12'b111111111111;
assign CPM[8128] = 12'b111111111111;
assign CPM[8129] = 12'b111111111111;
assign CPM[8130] = 12'b111111111111;
assign CPM[8131] = 12'b111111111111;
assign CPM[8132] = 12'b111111111111;
assign CPM[8133] = 12'b111111111111;
assign CPM[8134] = 12'b111111111111;
assign CPM[8135] = 12'b111111111111;
assign CPM[8136] = 12'b111111111111;
assign CPM[8137] = 12'b111111111111;
assign CPM[8138] = 12'b111111111111;
assign CPM[8139] = 12'b111111111111;
assign CPM[8140] = 12'b111111111111;
assign CPM[8141] = 12'b111111111111;
assign CPM[8142] = 12'b111111111111;
assign CPM[8143] = 12'b111111111111;
assign CPM[8144] = 12'b111111111111;
assign CPM[8145] = 12'b111111111111;
assign CPM[8146] = 12'b111111111111;
assign CPM[8147] = 12'b111111111111;
assign CPM[8148] = 12'b111111111111;
assign CPM[8149] = 12'b111111111111;
assign CPM[8150] = 12'b111111111111;
assign CPM[8151] = 12'b111111111111;
assign CPM[8152] = 12'b111111111111;
assign CPM[8153] = 12'b111111111111;
assign CPM[8154] = 12'b111111111111;
assign CPM[8155] = 12'b111111111111;
assign CPM[8156] = 12'b111111111111;
assign CPM[8157] = 12'b111111111111;
assign CPM[8158] = 12'b111111111111;
assign CPM[8159] = 12'b111111111111;
assign CPM[8160] = 12'b111111111111;
assign CPM[8161] = 12'b111111111111;
assign CPM[8162] = 12'b111111111111;
assign CPM[8163] = 12'b111111111111;
assign CPM[8164] = 12'b111111111111;
assign CPM[8165] = 12'b111111111111;
assign CPM[8166] = 12'b111111111111;
assign CPM[8167] = 12'b111111111111;
assign CPM[8168] = 12'b111111111111;
assign CPM[8169] = 12'b111111111111;
assign CPM[8170] = 12'b111111111111;
assign CPM[8171] = 12'b111111111111;
assign CPM[8172] = 12'b111111111111;
assign CPM[8173] = 12'b111111111111;
assign CPM[8174] = 12'b111111111111;
assign CPM[8175] = 12'b111111111111;
assign CPM[8176] = 12'b111111111111;
assign CPM[8177] = 12'b111111111111;
assign CPM[8178] = 12'b111111111111;
assign CPM[8179] = 12'b111111111111;
assign CPM[8180] = 12'b111111111111;
assign CPM[8181] = 12'b111111111111;
assign CPM[8182] = 12'b111111111111;
assign CPM[8183] = 12'b111111111111;
assign CPM[8184] = 12'b111111111111;
assign CPM[8185] = 12'b111111111111;
assign CPM[8186] = 12'b111111111111;
assign CPM[8187] = 12'b111111111111;
assign CPM[8188] = 12'b111111111111;
assign CPM[8189] = 12'b111111111111;
assign CPM[8190] = 12'b111111111111;
assign CPM[8191] = 12'b111111111111;
assign CPM[8192] = 12'b111111111111;
assign CPM[8193] = 12'b111111111111;
assign CPM[8194] = 12'b111111111111;
assign CPM[8195] = 12'b111111111111;
assign CPM[8196] = 12'b111111111111;
assign CPM[8197] = 12'b111111111111;
assign CPM[8198] = 12'b111111111111;
assign CPM[8199] = 12'b111111111111;
assign CPM[8200] = 12'b111111111111;
assign CPM[8201] = 12'b111111111111;
assign CPM[8202] = 12'b111111111111;
assign CPM[8203] = 12'b111111111111;
assign CPM[8204] = 12'b111111111111;
assign CPM[8205] = 12'b111111111111;
assign CPM[8206] = 12'b111111111111;
assign CPM[8207] = 12'b111111111111;
assign CPM[8208] = 12'b111111111111;
assign CPM[8209] = 12'b111111111111;
assign CPM[8210] = 12'b111111111111;
assign CPM[8211] = 12'b111111111111;
assign CPM[8212] = 12'b111111111111;
assign CPM[8213] = 12'b111111111111;
assign CPM[8214] = 12'b111111111111;
assign CPM[8215] = 12'b111111111111;
assign CPM[8216] = 12'b111111111111;
assign CPM[8217] = 12'b111111111111;
assign CPM[8218] = 12'b111111111111;
assign CPM[8219] = 12'b111111111111;
assign CPM[8220] = 12'b111111111111;
assign CPM[8221] = 12'b111111111111;
assign CPM[8222] = 12'b111111111111;
assign CPM[8223] = 12'b111111111111;
assign CPM[8224] = 12'b111111111111;
assign CPM[8225] = 12'b111111111111;
assign CPM[8226] = 12'b111111111111;
assign CPM[8227] = 12'b111111111111;
assign CPM[8228] = 12'b111111111111;
assign CPM[8229] = 12'b111111111111;
assign CPM[8230] = 12'b111111111111;
assign CPM[8231] = 12'b111111111111;
assign CPM[8232] = 12'b111111111111;
assign CPM[8233] = 12'b111111111111;
assign CPM[8234] = 12'b111111111111;
assign CPM[8235] = 12'b111111111111;
assign CPM[8236] = 12'b111111111111;
assign CPM[8237] = 12'b111111111111;
assign CPM[8238] = 12'b111111111111;
assign CPM[8239] = 12'b111111111111;
assign CPM[8240] = 12'b111111111111;
assign CPM[8241] = 12'b111111111111;
assign CPM[8242] = 12'b111111111111;
assign CPM[8243] = 12'b111111111111;
assign CPM[8244] = 12'b111111111111;
assign CPM[8245] = 12'b111111111111;
assign CPM[8246] = 12'b111111111111;
assign CPM[8247] = 12'b111111111111;
assign CPM[8248] = 12'b111111111111;
assign CPM[8249] = 12'b111111111111;
assign CPM[8250] = 12'b111111111111;
assign CPM[8251] = 12'b111111111111;
assign CPM[8252] = 12'b111111111111;
assign CPM[8253] = 12'b111111111111;
assign CPM[8254] = 12'b111111111111;
assign CPM[8255] = 12'b111111111111;
assign CPM[8256] = 12'b111111111111;
assign CPM[8257] = 12'b111111111111;
assign CPM[8258] = 12'b111111111111;
assign CPM[8259] = 12'b111111111111;
assign CPM[8260] = 12'b111111111111;
assign CPM[8261] = 12'b111111111111;
assign CPM[8262] = 12'b111111111111;
assign CPM[8263] = 12'b111111111111;
assign CPM[8264] = 12'b111111111111;
assign CPM[8265] = 12'b111111111111;
assign CPM[8266] = 12'b111111111111;
assign CPM[8267] = 12'b111111111111;
assign CPM[8268] = 12'b111111111111;
assign CPM[8269] = 12'b111111111111;
assign CPM[8270] = 12'b111111111111;
assign CPM[8271] = 12'b111111111111;
assign CPM[8272] = 12'b111111111111;
assign CPM[8273] = 12'b111111111111;
assign CPM[8274] = 12'b111111111111;
assign CPM[8275] = 12'b111111111111;
assign CPM[8276] = 12'b111111111111;
assign CPM[8277] = 12'b111111111111;
assign CPM[8278] = 12'b111111111111;
assign CPM[8279] = 12'b111111111111;
assign CPM[8280] = 12'b111111111111;
assign CPM[8281] = 12'b111111111111;
assign CPM[8282] = 12'b111111111111;
assign CPM[8283] = 12'b111111111111;
assign CPM[8284] = 12'b111111111111;
assign CPM[8285] = 12'b111111111111;
assign CPM[8286] = 12'b111111111111;
assign CPM[8287] = 12'b111111111111;
assign CPM[8288] = 12'b111111111111;
assign CPM[8289] = 12'b111111111111;
assign CPM[8290] = 12'b111111111111;
assign CPM[8291] = 12'b111111111111;
assign CPM[8292] = 12'b111111111111;
assign CPM[8293] = 12'b111111111111;
assign CPM[8294] = 12'b111111111111;
assign CPM[8295] = 12'b111111111111;
assign CPM[8296] = 12'b000000000000;
assign CPM[8297] = 12'b000000000000;
assign CPM[8298] = 12'b000000000000;
assign CPM[8299] = 12'b000000000000;
assign CPM[8300] = 12'b000000000000;
assign CPM[8301] = 12'b000000000000;
assign CPM[8302] = 12'b000000000000;
assign CPM[8303] = 12'b000000000000;
assign CPM[8304] = 12'b000000000000;
assign CPM[8305] = 12'b000000000000;
assign CPM[8306] = 12'b000000000000;
assign CPM[8307] = 12'b000000000000;
assign CPM[8308] = 12'b000000000000;
assign CPM[8309] = 12'b000000000000;
assign CPM[8310] = 12'b000000000000;
assign CPM[8311] = 12'b000000000000;
assign CPM[8312] = 12'b000000000000;
assign CPM[8313] = 12'b111111111111;
assign CPM[8314] = 12'b111111111111;
assign CPM[8315] = 12'b111111111111;
assign CPM[8316] = 12'b111111111111;
assign CPM[8317] = 12'b111111111111;
assign CPM[8318] = 12'b111111111111;
assign CPM[8319] = 12'b111111111111;
assign CPM[8320] = 12'b111111111111;
assign CPM[8321] = 12'b111111111111;
assign CPM[8322] = 12'b111111111111;
assign CPM[8323] = 12'b111111111111;
assign CPM[8324] = 12'b111111111111;
assign CPM[8325] = 12'b111111111111;
assign CPM[8326] = 12'b111111111111;
assign CPM[8327] = 12'b111111111111;
assign CPM[8328] = 12'b000000000000;
assign CPM[8329] = 12'b000000000000;
assign CPM[8330] = 12'b000000000000;
assign CPM[8331] = 12'b000000000000;
assign CPM[8332] = 12'b000000000000;
assign CPM[8333] = 12'b000000000000;
assign CPM[8334] = 12'b000000000000;
assign CPM[8335] = 12'b000000000000;
assign CPM[8336] = 12'b000000000000;
assign CPM[8337] = 12'b000000000000;
assign CPM[8338] = 12'b000000000000;
assign CPM[8339] = 12'b000000000000;
assign CPM[8340] = 12'b000000000000;
assign CPM[8341] = 12'b000000000000;
assign CPM[8342] = 12'b000000000000;
assign CPM[8343] = 12'b000000000000;
assign CPM[8344] = 12'b000000000000;
assign CPM[8345] = 12'b111111111111;
assign CPM[8346] = 12'b111111111111;
assign CPM[8347] = 12'b111111111111;
assign CPM[8348] = 12'b111111111111;
assign CPM[8349] = 12'b111111111111;
assign CPM[8350] = 12'b111111111111;
assign CPM[8351] = 12'b111111111111;
assign CPM[8352] = 12'b111111111111;
assign CPM[8353] = 12'b111111111111;
assign CPM[8354] = 12'b111111111111;
assign CPM[8355] = 12'b111111111111;
assign CPM[8356] = 12'b111111111111;
assign CPM[8357] = 12'b111111111111;
assign CPM[8358] = 12'b111111111111;
assign CPM[8359] = 12'b111111111111;
assign CPM[8360] = 12'b000000000000;
assign CPM[8361] = 12'b000000000000;
assign CPM[8362] = 12'b000000000000;
assign CPM[8363] = 12'b000000000000;
assign CPM[8364] = 12'b000000000000;
assign CPM[8365] = 12'b000000000000;
assign CPM[8366] = 12'b000000000000;
assign CPM[8367] = 12'b000000000000;
assign CPM[8368] = 12'b000000000000;
assign CPM[8369] = 12'b000000000000;
assign CPM[8370] = 12'b000000000000;
assign CPM[8371] = 12'b000000000000;
assign CPM[8372] = 12'b000000000000;
assign CPM[8373] = 12'b000000000000;
assign CPM[8374] = 12'b000000000000;
assign CPM[8375] = 12'b000000000000;
assign CPM[8376] = 12'b000000000000;
assign CPM[8377] = 12'b111111111111;
assign CPM[8378] = 12'b111111111111;
assign CPM[8379] = 12'b111111111111;
assign CPM[8380] = 12'b111111111111;
assign CPM[8381] = 12'b111111111111;
assign CPM[8382] = 12'b111111111111;
assign CPM[8383] = 12'b111111111111;
assign CPM[8384] = 12'b111111111111;
assign CPM[8385] = 12'b111111111111;
assign CPM[8386] = 12'b111111111111;
assign CPM[8387] = 12'b111111111111;
assign CPM[8388] = 12'b111111111111;
assign CPM[8389] = 12'b111111111111;
assign CPM[8390] = 12'b111111111111;
assign CPM[8391] = 12'b111111111111;
assign CPM[8392] = 12'b000000000000;
assign CPM[8393] = 12'b000000000000;
assign CPM[8394] = 12'b000000000000;
assign CPM[8395] = 12'b000000000000;
assign CPM[8396] = 12'b000000000000;
assign CPM[8397] = 12'b000000000000;
assign CPM[8398] = 12'b000000000000;
assign CPM[8399] = 12'b000000000000;
assign CPM[8400] = 12'b000000000000;
assign CPM[8401] = 12'b000000000000;
assign CPM[8402] = 12'b000000000000;
assign CPM[8403] = 12'b000000000000;
assign CPM[8404] = 12'b000000000000;
assign CPM[8405] = 12'b000000000000;
assign CPM[8406] = 12'b000000000000;
assign CPM[8407] = 12'b000000000000;
assign CPM[8408] = 12'b000000000000;
assign CPM[8409] = 12'b111111111111;
assign CPM[8410] = 12'b111111111111;
assign CPM[8411] = 12'b111111111111;
assign CPM[8412] = 12'b111111111111;
assign CPM[8413] = 12'b111111111111;
assign CPM[8414] = 12'b111111111111;
assign CPM[8415] = 12'b111111111111;
assign CPM[8416] = 12'b111111111111;
assign CPM[8417] = 12'b111111111111;
assign CPM[8418] = 12'b111111111111;
assign CPM[8419] = 12'b111111111111;
assign CPM[8420] = 12'b111111111111;
assign CPM[8421] = 12'b111111111111;
assign CPM[8422] = 12'b111111111111;
assign CPM[8423] = 12'b111111111111;
assign CPM[8424] = 12'b000000000000;
assign CPM[8425] = 12'b000000000000;
assign CPM[8426] = 12'b000000000000;
assign CPM[8427] = 12'b000000000000;
assign CPM[8428] = 12'b111111111111;
assign CPM[8429] = 12'b111111111111;
assign CPM[8430] = 12'b111111111111;
assign CPM[8431] = 12'b111111111111;
assign CPM[8432] = 12'b111111111111;
assign CPM[8433] = 12'b111111111111;
assign CPM[8434] = 12'b111111111111;
assign CPM[8435] = 12'b111111111111;
assign CPM[8436] = 12'b111111111111;
assign CPM[8437] = 12'b111111111111;
assign CPM[8438] = 12'b111111111111;
assign CPM[8439] = 12'b111111111111;
assign CPM[8440] = 12'b111111111111;
assign CPM[8441] = 12'b111111111111;
assign CPM[8442] = 12'b111111111111;
assign CPM[8443] = 12'b111111111111;
assign CPM[8444] = 12'b111111111111;
assign CPM[8445] = 12'b111111111111;
assign CPM[8446] = 12'b111111111111;
assign CPM[8447] = 12'b111111111111;
assign CPM[8448] = 12'b111111111111;
assign CPM[8449] = 12'b111111111111;
assign CPM[8450] = 12'b111111111111;
assign CPM[8451] = 12'b111111111111;
assign CPM[8452] = 12'b111111111111;
assign CPM[8453] = 12'b111111111111;
assign CPM[8454] = 12'b111111111111;
assign CPM[8455] = 12'b111111111111;
assign CPM[8456] = 12'b000000000000;
assign CPM[8457] = 12'b000000000000;
assign CPM[8458] = 12'b000000000000;
assign CPM[8459] = 12'b000000000000;
assign CPM[8460] = 12'b111111111111;
assign CPM[8461] = 12'b111111111111;
assign CPM[8462] = 12'b111111111111;
assign CPM[8463] = 12'b111111111111;
assign CPM[8464] = 12'b111111111111;
assign CPM[8465] = 12'b111111111111;
assign CPM[8466] = 12'b111111111111;
assign CPM[8467] = 12'b111111111111;
assign CPM[8468] = 12'b111111111111;
assign CPM[8469] = 12'b111111111111;
assign CPM[8470] = 12'b111111111111;
assign CPM[8471] = 12'b111111111111;
assign CPM[8472] = 12'b111111111111;
assign CPM[8473] = 12'b111111111111;
assign CPM[8474] = 12'b111111111111;
assign CPM[8475] = 12'b111111111111;
assign CPM[8476] = 12'b111111111111;
assign CPM[8477] = 12'b111111111111;
assign CPM[8478] = 12'b111111111111;
assign CPM[8479] = 12'b111111111111;
assign CPM[8480] = 12'b111111111111;
assign CPM[8481] = 12'b111111111111;
assign CPM[8482] = 12'b111111111111;
assign CPM[8483] = 12'b111111111111;
assign CPM[8484] = 12'b111111111111;
assign CPM[8485] = 12'b111111111111;
assign CPM[8486] = 12'b111111111111;
assign CPM[8487] = 12'b111111111111;
assign CPM[8488] = 12'b000000000000;
assign CPM[8489] = 12'b000000000000;
assign CPM[8490] = 12'b000000000000;
assign CPM[8491] = 12'b000000000000;
assign CPM[8492] = 12'b111111111111;
assign CPM[8493] = 12'b111111111111;
assign CPM[8494] = 12'b111111111111;
assign CPM[8495] = 12'b111111111111;
assign CPM[8496] = 12'b111111111111;
assign CPM[8497] = 12'b111111111111;
assign CPM[8498] = 12'b111111111111;
assign CPM[8499] = 12'b111111111111;
assign CPM[8500] = 12'b111111111111;
assign CPM[8501] = 12'b111111111111;
assign CPM[8502] = 12'b111111111111;
assign CPM[8503] = 12'b111111111111;
assign CPM[8504] = 12'b111111111111;
assign CPM[8505] = 12'b111111111111;
assign CPM[8506] = 12'b111111111111;
assign CPM[8507] = 12'b111111111111;
assign CPM[8508] = 12'b111111111111;
assign CPM[8509] = 12'b111111111111;
assign CPM[8510] = 12'b111111111111;
assign CPM[8511] = 12'b111111111111;
assign CPM[8512] = 12'b111111111111;
assign CPM[8513] = 12'b111111111111;
assign CPM[8514] = 12'b111111111111;
assign CPM[8515] = 12'b111111111111;
assign CPM[8516] = 12'b111111111111;
assign CPM[8517] = 12'b111111111111;
assign CPM[8518] = 12'b111111111111;
assign CPM[8519] = 12'b111111111111;
assign CPM[8520] = 12'b000000000000;
assign CPM[8521] = 12'b000000000000;
assign CPM[8522] = 12'b000000000000;
assign CPM[8523] = 12'b000000000000;
assign CPM[8524] = 12'b111111111111;
assign CPM[8525] = 12'b111111111111;
assign CPM[8526] = 12'b111111111111;
assign CPM[8527] = 12'b111111111111;
assign CPM[8528] = 12'b111111111111;
assign CPM[8529] = 12'b111111111111;
assign CPM[8530] = 12'b111111111111;
assign CPM[8531] = 12'b111111111111;
assign CPM[8532] = 12'b111111111111;
assign CPM[8533] = 12'b111111111111;
assign CPM[8534] = 12'b111111111111;
assign CPM[8535] = 12'b111111111111;
assign CPM[8536] = 12'b111111111111;
assign CPM[8537] = 12'b111111111111;
assign CPM[8538] = 12'b111111111111;
assign CPM[8539] = 12'b111111111111;
assign CPM[8540] = 12'b111111111111;
assign CPM[8541] = 12'b111111111111;
assign CPM[8542] = 12'b111111111111;
assign CPM[8543] = 12'b111111111111;
assign CPM[8544] = 12'b111111111111;
assign CPM[8545] = 12'b111111111111;
assign CPM[8546] = 12'b111111111111;
assign CPM[8547] = 12'b111111111111;
assign CPM[8548] = 12'b111111111111;
assign CPM[8549] = 12'b111111111111;
assign CPM[8550] = 12'b111111111111;
assign CPM[8551] = 12'b111111111111;
assign CPM[8552] = 12'b000000000000;
assign CPM[8553] = 12'b000000000000;
assign CPM[8554] = 12'b000000000000;
assign CPM[8555] = 12'b000000000000;
assign CPM[8556] = 12'b111111111111;
assign CPM[8557] = 12'b111111111111;
assign CPM[8558] = 12'b111111111111;
assign CPM[8559] = 12'b111111111111;
assign CPM[8560] = 12'b111111111111;
assign CPM[8561] = 12'b111111111111;
assign CPM[8562] = 12'b111111111111;
assign CPM[8563] = 12'b111111111111;
assign CPM[8564] = 12'b111111111111;
assign CPM[8565] = 12'b111111111111;
assign CPM[8566] = 12'b111111111111;
assign CPM[8567] = 12'b111111111111;
assign CPM[8568] = 12'b111111111111;
assign CPM[8569] = 12'b111111111111;
assign CPM[8570] = 12'b111111111111;
assign CPM[8571] = 12'b111111111111;
assign CPM[8572] = 12'b111111111111;
assign CPM[8573] = 12'b111111111111;
assign CPM[8574] = 12'b111111111111;
assign CPM[8575] = 12'b111111111111;
assign CPM[8576] = 12'b111111111111;
assign CPM[8577] = 12'b111111111111;
assign CPM[8578] = 12'b111111111111;
assign CPM[8579] = 12'b111111111111;
assign CPM[8580] = 12'b111111111111;
assign CPM[8581] = 12'b111111111111;
assign CPM[8582] = 12'b111111111111;
assign CPM[8583] = 12'b111111111111;
assign CPM[8584] = 12'b000000000000;
assign CPM[8585] = 12'b000000000000;
assign CPM[8586] = 12'b000000000000;
assign CPM[8587] = 12'b000000000000;
assign CPM[8588] = 12'b111111111111;
assign CPM[8589] = 12'b111111111111;
assign CPM[8590] = 12'b111111111111;
assign CPM[8591] = 12'b111111111111;
assign CPM[8592] = 12'b111111111111;
assign CPM[8593] = 12'b111111111111;
assign CPM[8594] = 12'b111111111111;
assign CPM[8595] = 12'b111111111111;
assign CPM[8596] = 12'b111111111111;
assign CPM[8597] = 12'b111111111111;
assign CPM[8598] = 12'b111111111111;
assign CPM[8599] = 12'b111111111111;
assign CPM[8600] = 12'b111111111111;
assign CPM[8601] = 12'b111111111111;
assign CPM[8602] = 12'b111111111111;
assign CPM[8603] = 12'b111111111111;
assign CPM[8604] = 12'b111111111111;
assign CPM[8605] = 12'b111111111111;
assign CPM[8606] = 12'b111111111111;
assign CPM[8607] = 12'b111111111111;
assign CPM[8608] = 12'b111111111111;
assign CPM[8609] = 12'b111111111111;
assign CPM[8610] = 12'b111111111111;
assign CPM[8611] = 12'b111111111111;
assign CPM[8612] = 12'b111111111111;
assign CPM[8613] = 12'b111111111111;
assign CPM[8614] = 12'b111111111111;
assign CPM[8615] = 12'b111111111111;
assign CPM[8616] = 12'b000000000000;
assign CPM[8617] = 12'b000000000000;
assign CPM[8618] = 12'b000000000000;
assign CPM[8619] = 12'b000000000000;
assign CPM[8620] = 12'b111111111111;
assign CPM[8621] = 12'b111111111111;
assign CPM[8622] = 12'b111111111111;
assign CPM[8623] = 12'b111111111111;
assign CPM[8624] = 12'b111111111111;
assign CPM[8625] = 12'b111111111111;
assign CPM[8626] = 12'b111111111111;
assign CPM[8627] = 12'b111111111111;
assign CPM[8628] = 12'b111111111111;
assign CPM[8629] = 12'b111111111111;
assign CPM[8630] = 12'b111111111111;
assign CPM[8631] = 12'b111111111111;
assign CPM[8632] = 12'b111111111111;
assign CPM[8633] = 12'b111111111111;
assign CPM[8634] = 12'b111111111111;
assign CPM[8635] = 12'b111111111111;
assign CPM[8636] = 12'b111111111111;
assign CPM[8637] = 12'b111111111111;
assign CPM[8638] = 12'b111111111111;
assign CPM[8639] = 12'b111111111111;
assign CPM[8640] = 12'b111111111111;
assign CPM[8641] = 12'b111111111111;
assign CPM[8642] = 12'b111111111111;
assign CPM[8643] = 12'b111111111111;
assign CPM[8644] = 12'b111111111111;
assign CPM[8645] = 12'b111111111111;
assign CPM[8646] = 12'b111111111111;
assign CPM[8647] = 12'b111111111111;
assign CPM[8648] = 12'b000000000000;
assign CPM[8649] = 12'b000000000000;
assign CPM[8650] = 12'b000000000000;
assign CPM[8651] = 12'b000000000000;
assign CPM[8652] = 12'b111111111111;
assign CPM[8653] = 12'b111111111111;
assign CPM[8654] = 12'b111111111111;
assign CPM[8655] = 12'b111111111111;
assign CPM[8656] = 12'b111111111111;
assign CPM[8657] = 12'b111111111111;
assign CPM[8658] = 12'b111111111111;
assign CPM[8659] = 12'b111111111111;
assign CPM[8660] = 12'b111111111111;
assign CPM[8661] = 12'b111111111111;
assign CPM[8662] = 12'b111111111111;
assign CPM[8663] = 12'b111111111111;
assign CPM[8664] = 12'b111111111111;
assign CPM[8665] = 12'b111111111111;
assign CPM[8666] = 12'b111111111111;
assign CPM[8667] = 12'b111111111111;
assign CPM[8668] = 12'b111111111111;
assign CPM[8669] = 12'b111111111111;
assign CPM[8670] = 12'b111111111111;
assign CPM[8671] = 12'b111111111111;
assign CPM[8672] = 12'b111111111111;
assign CPM[8673] = 12'b111111111111;
assign CPM[8674] = 12'b111111111111;
assign CPM[8675] = 12'b111111111111;
assign CPM[8676] = 12'b111111111111;
assign CPM[8677] = 12'b111111111111;
assign CPM[8678] = 12'b111111111111;
assign CPM[8679] = 12'b111111111111;
assign CPM[8680] = 12'b111111111111;
assign CPM[8681] = 12'b111111111111;
assign CPM[8682] = 12'b111111111111;
assign CPM[8683] = 12'b111111111111;
assign CPM[8684] = 12'b000000000000;
assign CPM[8685] = 12'b000000000000;
assign CPM[8686] = 12'b000000000000;
assign CPM[8687] = 12'b000000000000;
assign CPM[8688] = 12'b000000000000;
assign CPM[8689] = 12'b000000000000;
assign CPM[8690] = 12'b000000000000;
assign CPM[8691] = 12'b000000000000;
assign CPM[8692] = 12'b000000000000;
assign CPM[8693] = 12'b000000000000;
assign CPM[8694] = 12'b000000000000;
assign CPM[8695] = 12'b111111111111;
assign CPM[8696] = 12'b111111111111;
assign CPM[8697] = 12'b111111111111;
assign CPM[8698] = 12'b111111111111;
assign CPM[8699] = 12'b111111111111;
assign CPM[8700] = 12'b111111111111;
assign CPM[8701] = 12'b111111111111;
assign CPM[8702] = 12'b111111111111;
assign CPM[8703] = 12'b111111111111;
assign CPM[8704] = 12'b111111111111;
assign CPM[8705] = 12'b111111111111;
assign CPM[8706] = 12'b111111111111;
assign CPM[8707] = 12'b111111111111;
assign CPM[8708] = 12'b111111111111;
assign CPM[8709] = 12'b111111111111;
assign CPM[8710] = 12'b111111111111;
assign CPM[8711] = 12'b111111111111;
assign CPM[8712] = 12'b111111111111;
assign CPM[8713] = 12'b111111111111;
assign CPM[8714] = 12'b111111111111;
assign CPM[8715] = 12'b111111111111;
assign CPM[8716] = 12'b000000000000;
assign CPM[8717] = 12'b000000000000;
assign CPM[8718] = 12'b000000000000;
assign CPM[8719] = 12'b000000000000;
assign CPM[8720] = 12'b000000000000;
assign CPM[8721] = 12'b000000000000;
assign CPM[8722] = 12'b000000000000;
assign CPM[8723] = 12'b000000000000;
assign CPM[8724] = 12'b000000000000;
assign CPM[8725] = 12'b000000000000;
assign CPM[8726] = 12'b000000000000;
assign CPM[8727] = 12'b111111111111;
assign CPM[8728] = 12'b111111111111;
assign CPM[8729] = 12'b111111111111;
assign CPM[8730] = 12'b111111111111;
assign CPM[8731] = 12'b111111111111;
assign CPM[8732] = 12'b111111111111;
assign CPM[8733] = 12'b111111111111;
assign CPM[8734] = 12'b111111111111;
assign CPM[8735] = 12'b111111111111;
assign CPM[8736] = 12'b111111111111;
assign CPM[8737] = 12'b111111111111;
assign CPM[8738] = 12'b111111111111;
assign CPM[8739] = 12'b111111111111;
assign CPM[8740] = 12'b111111111111;
assign CPM[8741] = 12'b111111111111;
assign CPM[8742] = 12'b111111111111;
assign CPM[8743] = 12'b111111111111;
assign CPM[8744] = 12'b111111111111;
assign CPM[8745] = 12'b111111111111;
assign CPM[8746] = 12'b111111111111;
assign CPM[8747] = 12'b111111111111;
assign CPM[8748] = 12'b000000000000;
assign CPM[8749] = 12'b000000000000;
assign CPM[8750] = 12'b000000000000;
assign CPM[8751] = 12'b000000000000;
assign CPM[8752] = 12'b000000000000;
assign CPM[8753] = 12'b000000000000;
assign CPM[8754] = 12'b000000000000;
assign CPM[8755] = 12'b000000000000;
assign CPM[8756] = 12'b000000000000;
assign CPM[8757] = 12'b000000000000;
assign CPM[8758] = 12'b000000000000;
assign CPM[8759] = 12'b111111111111;
assign CPM[8760] = 12'b111111111111;
assign CPM[8761] = 12'b111111111111;
assign CPM[8762] = 12'b111111111111;
assign CPM[8763] = 12'b111111111111;
assign CPM[8764] = 12'b111111111111;
assign CPM[8765] = 12'b111111111111;
assign CPM[8766] = 12'b111111111111;
assign CPM[8767] = 12'b111111111111;
assign CPM[8768] = 12'b111111111111;
assign CPM[8769] = 12'b111111111111;
assign CPM[8770] = 12'b111111111111;
assign CPM[8771] = 12'b111111111111;
assign CPM[8772] = 12'b111111111111;
assign CPM[8773] = 12'b111111111111;
assign CPM[8774] = 12'b111111111111;
assign CPM[8775] = 12'b111111111111;
assign CPM[8776] = 12'b111111111111;
assign CPM[8777] = 12'b111111111111;
assign CPM[8778] = 12'b111111111111;
assign CPM[8779] = 12'b111111111111;
assign CPM[8780] = 12'b000000000000;
assign CPM[8781] = 12'b000000000000;
assign CPM[8782] = 12'b000000000000;
assign CPM[8783] = 12'b000000000000;
assign CPM[8784] = 12'b000000000000;
assign CPM[8785] = 12'b000000000000;
assign CPM[8786] = 12'b000000000000;
assign CPM[8787] = 12'b000000000000;
assign CPM[8788] = 12'b000000000000;
assign CPM[8789] = 12'b000000000000;
assign CPM[8790] = 12'b000000000000;
assign CPM[8791] = 12'b111111111111;
assign CPM[8792] = 12'b111111111111;
assign CPM[8793] = 12'b111111111111;
assign CPM[8794] = 12'b111111111111;
assign CPM[8795] = 12'b111111111111;
assign CPM[8796] = 12'b111111111111;
assign CPM[8797] = 12'b111111111111;
assign CPM[8798] = 12'b111111111111;
assign CPM[8799] = 12'b111111111111;
assign CPM[8800] = 12'b111111111111;
assign CPM[8801] = 12'b111111111111;
assign CPM[8802] = 12'b111111111111;
assign CPM[8803] = 12'b111111111111;
assign CPM[8804] = 12'b111111111111;
assign CPM[8805] = 12'b111111111111;
assign CPM[8806] = 12'b111111111111;
assign CPM[8807] = 12'b111111111111;
assign CPM[8808] = 12'b111111111111;
assign CPM[8809] = 12'b111111111111;
assign CPM[8810] = 12'b111111111111;
assign CPM[8811] = 12'b111111111111;
assign CPM[8812] = 12'b111111111111;
assign CPM[8813] = 12'b111111111111;
assign CPM[8814] = 12'b111111111111;
assign CPM[8815] = 12'b111111111111;
assign CPM[8816] = 12'b111111111111;
assign CPM[8817] = 12'b111111111111;
assign CPM[8818] = 12'b111111111111;
assign CPM[8819] = 12'b111111111111;
assign CPM[8820] = 12'b111111111111;
assign CPM[8821] = 12'b111111111111;
assign CPM[8822] = 12'b111111111111;
assign CPM[8823] = 12'b000000000000;
assign CPM[8824] = 12'b000000000000;
assign CPM[8825] = 12'b000000000000;
assign CPM[8826] = 12'b000000000000;
assign CPM[8827] = 12'b111111111111;
assign CPM[8828] = 12'b111111111111;
assign CPM[8829] = 12'b111111111111;
assign CPM[8830] = 12'b111111111111;
assign CPM[8831] = 12'b111111111111;
assign CPM[8832] = 12'b111111111111;
assign CPM[8833] = 12'b111111111111;
assign CPM[8834] = 12'b111111111111;
assign CPM[8835] = 12'b111111111111;
assign CPM[8836] = 12'b111111111111;
assign CPM[8837] = 12'b111111111111;
assign CPM[8838] = 12'b111111111111;
assign CPM[8839] = 12'b111111111111;
assign CPM[8840] = 12'b111111111111;
assign CPM[8841] = 12'b111111111111;
assign CPM[8842] = 12'b111111111111;
assign CPM[8843] = 12'b111111111111;
assign CPM[8844] = 12'b111111111111;
assign CPM[8845] = 12'b111111111111;
assign CPM[8846] = 12'b111111111111;
assign CPM[8847] = 12'b111111111111;
assign CPM[8848] = 12'b111111111111;
assign CPM[8849] = 12'b111111111111;
assign CPM[8850] = 12'b111111111111;
assign CPM[8851] = 12'b111111111111;
assign CPM[8852] = 12'b111111111111;
assign CPM[8853] = 12'b111111111111;
assign CPM[8854] = 12'b111111111111;
assign CPM[8855] = 12'b000000000000;
assign CPM[8856] = 12'b000000000000;
assign CPM[8857] = 12'b000000000000;
assign CPM[8858] = 12'b000000000000;
assign CPM[8859] = 12'b111111111111;
assign CPM[8860] = 12'b111111111111;
assign CPM[8861] = 12'b111111111111;
assign CPM[8862] = 12'b111111111111;
assign CPM[8863] = 12'b111111111111;
assign CPM[8864] = 12'b111111111111;
assign CPM[8865] = 12'b111111111111;
assign CPM[8866] = 12'b111111111111;
assign CPM[8867] = 12'b111111111111;
assign CPM[8868] = 12'b111111111111;
assign CPM[8869] = 12'b111111111111;
assign CPM[8870] = 12'b111111111111;
assign CPM[8871] = 12'b111111111111;
assign CPM[8872] = 12'b111111111111;
assign CPM[8873] = 12'b111111111111;
assign CPM[8874] = 12'b111111111111;
assign CPM[8875] = 12'b111111111111;
assign CPM[8876] = 12'b111111111111;
assign CPM[8877] = 12'b111111111111;
assign CPM[8878] = 12'b111111111111;
assign CPM[8879] = 12'b111111111111;
assign CPM[8880] = 12'b111111111111;
assign CPM[8881] = 12'b111111111111;
assign CPM[8882] = 12'b111111111111;
assign CPM[8883] = 12'b111111111111;
assign CPM[8884] = 12'b111111111111;
assign CPM[8885] = 12'b111111111111;
assign CPM[8886] = 12'b111111111111;
assign CPM[8887] = 12'b000000000000;
assign CPM[8888] = 12'b000000000000;
assign CPM[8889] = 12'b000000000000;
assign CPM[8890] = 12'b000000000000;
assign CPM[8891] = 12'b111111111111;
assign CPM[8892] = 12'b111111111111;
assign CPM[8893] = 12'b111111111111;
assign CPM[8894] = 12'b111111111111;
assign CPM[8895] = 12'b111111111111;
assign CPM[8896] = 12'b111111111111;
assign CPM[8897] = 12'b111111111111;
assign CPM[8898] = 12'b111111111111;
assign CPM[8899] = 12'b111111111111;
assign CPM[8900] = 12'b111111111111;
assign CPM[8901] = 12'b111111111111;
assign CPM[8902] = 12'b111111111111;
assign CPM[8903] = 12'b111111111111;
assign CPM[8904] = 12'b111111111111;
assign CPM[8905] = 12'b111111111111;
assign CPM[8906] = 12'b111111111111;
assign CPM[8907] = 12'b111111111111;
assign CPM[8908] = 12'b111111111111;
assign CPM[8909] = 12'b111111111111;
assign CPM[8910] = 12'b111111111111;
assign CPM[8911] = 12'b111111111111;
assign CPM[8912] = 12'b111111111111;
assign CPM[8913] = 12'b111111111111;
assign CPM[8914] = 12'b111111111111;
assign CPM[8915] = 12'b111111111111;
assign CPM[8916] = 12'b111111111111;
assign CPM[8917] = 12'b111111111111;
assign CPM[8918] = 12'b111111111111;
assign CPM[8919] = 12'b000000000000;
assign CPM[8920] = 12'b000000000000;
assign CPM[8921] = 12'b000000000000;
assign CPM[8922] = 12'b000000000000;
assign CPM[8923] = 12'b111111111111;
assign CPM[8924] = 12'b111111111111;
assign CPM[8925] = 12'b111111111111;
assign CPM[8926] = 12'b111111111111;
assign CPM[8927] = 12'b111111111111;
assign CPM[8928] = 12'b111111111111;
assign CPM[8929] = 12'b111111111111;
assign CPM[8930] = 12'b111111111111;
assign CPM[8931] = 12'b111111111111;
assign CPM[8932] = 12'b111111111111;
assign CPM[8933] = 12'b111111111111;
assign CPM[8934] = 12'b000000000000;
assign CPM[8935] = 12'b000000000000;
assign CPM[8936] = 12'b000000000000;
assign CPM[8937] = 12'b000000000000;
assign CPM[8938] = 12'b111111111111;
assign CPM[8939] = 12'b111111111111;
assign CPM[8940] = 12'b111111111111;
assign CPM[8941] = 12'b111111111111;
assign CPM[8942] = 12'b111111111111;
assign CPM[8943] = 12'b111111111111;
assign CPM[8944] = 12'b111111111111;
assign CPM[8945] = 12'b111111111111;
assign CPM[8946] = 12'b111111111111;
assign CPM[8947] = 12'b111111111111;
assign CPM[8948] = 12'b111111111111;
assign CPM[8949] = 12'b111111111111;
assign CPM[8950] = 12'b111111111111;
assign CPM[8951] = 12'b000000000000;
assign CPM[8952] = 12'b000000000000;
assign CPM[8953] = 12'b000000000000;
assign CPM[8954] = 12'b000000000000;
assign CPM[8955] = 12'b111111111111;
assign CPM[8956] = 12'b111111111111;
assign CPM[8957] = 12'b111111111111;
assign CPM[8958] = 12'b111111111111;
assign CPM[8959] = 12'b111111111111;
assign CPM[8960] = 12'b111111111111;
assign CPM[8961] = 12'b111111111111;
assign CPM[8962] = 12'b111111111111;
assign CPM[8963] = 12'b111111111111;
assign CPM[8964] = 12'b111111111111;
assign CPM[8965] = 12'b111111111111;
assign CPM[8966] = 12'b000000000000;
assign CPM[8967] = 12'b000000000000;
assign CPM[8968] = 12'b000000000000;
assign CPM[8969] = 12'b000000000000;
assign CPM[8970] = 12'b111111111111;
assign CPM[8971] = 12'b111111111111;
assign CPM[8972] = 12'b111111111111;
assign CPM[8973] = 12'b111111111111;
assign CPM[8974] = 12'b111111111111;
assign CPM[8975] = 12'b111111111111;
assign CPM[8976] = 12'b111111111111;
assign CPM[8977] = 12'b111111111111;
assign CPM[8978] = 12'b111111111111;
assign CPM[8979] = 12'b111111111111;
assign CPM[8980] = 12'b111111111111;
assign CPM[8981] = 12'b111111111111;
assign CPM[8982] = 12'b111111111111;
assign CPM[8983] = 12'b000000000000;
assign CPM[8984] = 12'b000000000000;
assign CPM[8985] = 12'b000000000000;
assign CPM[8986] = 12'b000000000000;
assign CPM[8987] = 12'b111111111111;
assign CPM[8988] = 12'b111111111111;
assign CPM[8989] = 12'b111111111111;
assign CPM[8990] = 12'b111111111111;
assign CPM[8991] = 12'b111111111111;
assign CPM[8992] = 12'b111111111111;
assign CPM[8993] = 12'b111111111111;
assign CPM[8994] = 12'b111111111111;
assign CPM[8995] = 12'b111111111111;
assign CPM[8996] = 12'b111111111111;
assign CPM[8997] = 12'b111111111111;
assign CPM[8998] = 12'b000000000000;
assign CPM[8999] = 12'b000000000000;
assign CPM[9000] = 12'b000000000000;
assign CPM[9001] = 12'b000000000000;
assign CPM[9002] = 12'b111111111111;
assign CPM[9003] = 12'b111111111111;
assign CPM[9004] = 12'b111111111111;
assign CPM[9005] = 12'b111111111111;
assign CPM[9006] = 12'b111111111111;
assign CPM[9007] = 12'b111111111111;
assign CPM[9008] = 12'b111111111111;
assign CPM[9009] = 12'b111111111111;
assign CPM[9010] = 12'b111111111111;
assign CPM[9011] = 12'b111111111111;
assign CPM[9012] = 12'b111111111111;
assign CPM[9013] = 12'b111111111111;
assign CPM[9014] = 12'b111111111111;
assign CPM[9015] = 12'b000000000000;
assign CPM[9016] = 12'b000000000000;
assign CPM[9017] = 12'b000000000000;
assign CPM[9018] = 12'b000000000000;
assign CPM[9019] = 12'b111111111111;
assign CPM[9020] = 12'b111111111111;
assign CPM[9021] = 12'b111111111111;
assign CPM[9022] = 12'b111111111111;
assign CPM[9023] = 12'b111111111111;
assign CPM[9024] = 12'b111111111111;
assign CPM[9025] = 12'b111111111111;
assign CPM[9026] = 12'b111111111111;
assign CPM[9027] = 12'b111111111111;
assign CPM[9028] = 12'b111111111111;
assign CPM[9029] = 12'b111111111111;
assign CPM[9030] = 12'b000000000000;
assign CPM[9031] = 12'b000000000000;
assign CPM[9032] = 12'b000000000000;
assign CPM[9033] = 12'b000000000000;
assign CPM[9034] = 12'b111111111111;
assign CPM[9035] = 12'b111111111111;
assign CPM[9036] = 12'b111111111111;
assign CPM[9037] = 12'b111111111111;
assign CPM[9038] = 12'b111111111111;
assign CPM[9039] = 12'b111111111111;
assign CPM[9040] = 12'b111111111111;
assign CPM[9041] = 12'b111111111111;
assign CPM[9042] = 12'b111111111111;
assign CPM[9043] = 12'b111111111111;
assign CPM[9044] = 12'b111111111111;
assign CPM[9045] = 12'b111111111111;
assign CPM[9046] = 12'b111111111111;
assign CPM[9047] = 12'b000000000000;
assign CPM[9048] = 12'b000000000000;
assign CPM[9049] = 12'b000000000000;
assign CPM[9050] = 12'b000000000000;
assign CPM[9051] = 12'b111111111111;
assign CPM[9052] = 12'b111111111111;
assign CPM[9053] = 12'b111111111111;
assign CPM[9054] = 12'b111111111111;
assign CPM[9055] = 12'b111111111111;
assign CPM[9056] = 12'b111111111111;
assign CPM[9057] = 12'b111111111111;
assign CPM[9058] = 12'b111111111111;
assign CPM[9059] = 12'b111111111111;
assign CPM[9060] = 12'b111111111111;
assign CPM[9061] = 12'b111111111111;
assign CPM[9062] = 12'b111111111111;
assign CPM[9063] = 12'b111111111111;
assign CPM[9064] = 12'b111111111111;
assign CPM[9065] = 12'b111111111111;
assign CPM[9066] = 12'b000000000000;
assign CPM[9067] = 12'b000000000000;
assign CPM[9068] = 12'b000000000000;
assign CPM[9069] = 12'b000000000000;
assign CPM[9070] = 12'b000000000000;
assign CPM[9071] = 12'b000000000000;
assign CPM[9072] = 12'b000000000000;
assign CPM[9073] = 12'b000000000000;
assign CPM[9074] = 12'b000000000000;
assign CPM[9075] = 12'b000000000000;
assign CPM[9076] = 12'b000000000000;
assign CPM[9077] = 12'b000000000000;
assign CPM[9078] = 12'b000000000000;
assign CPM[9079] = 12'b111111111111;
assign CPM[9080] = 12'b111111111111;
assign CPM[9081] = 12'b111111111111;
assign CPM[9082] = 12'b111111111111;
assign CPM[9083] = 12'b111111111111;
assign CPM[9084] = 12'b111111111111;
assign CPM[9085] = 12'b111111111111;
assign CPM[9086] = 12'b111111111111;
assign CPM[9087] = 12'b111111111111;
assign CPM[9088] = 12'b111111111111;
assign CPM[9089] = 12'b111111111111;
assign CPM[9090] = 12'b111111111111;
assign CPM[9091] = 12'b111111111111;
assign CPM[9092] = 12'b111111111111;
assign CPM[9093] = 12'b111111111111;
assign CPM[9094] = 12'b111111111111;
assign CPM[9095] = 12'b111111111111;
assign CPM[9096] = 12'b111111111111;
assign CPM[9097] = 12'b111111111111;
assign CPM[9098] = 12'b000000000000;
assign CPM[9099] = 12'b000000000000;
assign CPM[9100] = 12'b000000000000;
assign CPM[9101] = 12'b000000000000;
assign CPM[9102] = 12'b000000000000;
assign CPM[9103] = 12'b000000000000;
assign CPM[9104] = 12'b000000000000;
assign CPM[9105] = 12'b000000000000;
assign CPM[9106] = 12'b000000000000;
assign CPM[9107] = 12'b000000000000;
assign CPM[9108] = 12'b000000000000;
assign CPM[9109] = 12'b000000000000;
assign CPM[9110] = 12'b000000000000;
assign CPM[9111] = 12'b111111111111;
assign CPM[9112] = 12'b111111111111;
assign CPM[9113] = 12'b111111111111;
assign CPM[9114] = 12'b111111111111;
assign CPM[9115] = 12'b111111111111;
assign CPM[9116] = 12'b111111111111;
assign CPM[9117] = 12'b111111111111;
assign CPM[9118] = 12'b111111111111;
assign CPM[9119] = 12'b111111111111;
assign CPM[9120] = 12'b111111111111;
assign CPM[9121] = 12'b111111111111;
assign CPM[9122] = 12'b111111111111;
assign CPM[9123] = 12'b111111111111;
assign CPM[9124] = 12'b111111111111;
assign CPM[9125] = 12'b111111111111;
assign CPM[9126] = 12'b111111111111;
assign CPM[9127] = 12'b111111111111;
assign CPM[9128] = 12'b111111111111;
assign CPM[9129] = 12'b111111111111;
assign CPM[9130] = 12'b000000000000;
assign CPM[9131] = 12'b000000000000;
assign CPM[9132] = 12'b000000000000;
assign CPM[9133] = 12'b000000000000;
assign CPM[9134] = 12'b000000000000;
assign CPM[9135] = 12'b000000000000;
assign CPM[9136] = 12'b000000000000;
assign CPM[9137] = 12'b000000000000;
assign CPM[9138] = 12'b000000000000;
assign CPM[9139] = 12'b000000000000;
assign CPM[9140] = 12'b000000000000;
assign CPM[9141] = 12'b000000000000;
assign CPM[9142] = 12'b000000000000;
assign CPM[9143] = 12'b111111111111;
assign CPM[9144] = 12'b111111111111;
assign CPM[9145] = 12'b111111111111;
assign CPM[9146] = 12'b111111111111;
assign CPM[9147] = 12'b111111111111;
assign CPM[9148] = 12'b111111111111;
assign CPM[9149] = 12'b111111111111;
assign CPM[9150] = 12'b111111111111;
assign CPM[9151] = 12'b111111111111;
assign CPM[9152] = 12'b111111111111;
assign CPM[9153] = 12'b111111111111;
assign CPM[9154] = 12'b111111111111;
assign CPM[9155] = 12'b111111111111;
assign CPM[9156] = 12'b111111111111;
assign CPM[9157] = 12'b111111111111;
assign CPM[9158] = 12'b111111111111;
assign CPM[9159] = 12'b111111111111;
assign CPM[9160] = 12'b111111111111;
assign CPM[9161] = 12'b111111111111;
assign CPM[9162] = 12'b000000000000;
assign CPM[9163] = 12'b000000000000;
assign CPM[9164] = 12'b000000000000;
assign CPM[9165] = 12'b000000000000;
assign CPM[9166] = 12'b000000000000;
assign CPM[9167] = 12'b000000000000;
assign CPM[9168] = 12'b000000000000;
assign CPM[9169] = 12'b000000000000;
assign CPM[9170] = 12'b000000000000;
assign CPM[9171] = 12'b000000000000;
assign CPM[9172] = 12'b000000000000;
assign CPM[9173] = 12'b000000000000;
assign CPM[9174] = 12'b000000000000;
assign CPM[9175] = 12'b111111111111;
assign CPM[9176] = 12'b111111111111;
assign CPM[9177] = 12'b111111111111;
assign CPM[9178] = 12'b111111111111;
assign CPM[9179] = 12'b111111111111;
assign CPM[9180] = 12'b111111111111;
assign CPM[9181] = 12'b111111111111;
assign CPM[9182] = 12'b111111111111;
assign CPM[9183] = 12'b111111111111;
assign CPM[9184] = 12'b111111111111;
assign CPM[9185] = 12'b111111111111;
assign CPM[9186] = 12'b111111111111;
assign CPM[9187] = 12'b111111111111;
assign CPM[9188] = 12'b111111111111;
assign CPM[9189] = 12'b111111111111;
assign CPM[9190] = 12'b111111111111;
assign CPM[9191] = 12'b111111111111;
assign CPM[9192] = 12'b111111111111;
assign CPM[9193] = 12'b111111111111;
assign CPM[9194] = 12'b111111111111;
assign CPM[9195] = 12'b111111111111;
assign CPM[9196] = 12'b111111111111;
assign CPM[9197] = 12'b111111111111;
assign CPM[9198] = 12'b111111111111;
assign CPM[9199] = 12'b111111111111;
assign CPM[9200] = 12'b111111111111;
assign CPM[9201] = 12'b111111111111;
assign CPM[9202] = 12'b111111111111;
assign CPM[9203] = 12'b111111111111;
assign CPM[9204] = 12'b111111111111;
assign CPM[9205] = 12'b111111111111;
assign CPM[9206] = 12'b111111111111;
assign CPM[9207] = 12'b111111111111;
assign CPM[9208] = 12'b111111111111;
assign CPM[9209] = 12'b111111111111;
assign CPM[9210] = 12'b111111111111;
assign CPM[9211] = 12'b111111111111;
assign CPM[9212] = 12'b111111111111;
assign CPM[9213] = 12'b111111111111;
assign CPM[9214] = 12'b111111111111;
assign CPM[9215] = 12'b111111111111;
assign CPM[9216] = 12'b111111111111;
assign CPM[9217] = 12'b111111111111;
assign CPM[9218] = 12'b111111111111;
assign CPM[9219] = 12'b111111111111;
assign CPM[9220] = 12'b111111111111;
assign CPM[9221] = 12'b111111111111;
assign CPM[9222] = 12'b111111111111;
assign CPM[9223] = 12'b111111111111;
assign CPM[9224] = 12'b111111111111;
assign CPM[9225] = 12'b111111111111;
assign CPM[9226] = 12'b111111111111;
assign CPM[9227] = 12'b111111111111;
assign CPM[9228] = 12'b111111111111;
assign CPM[9229] = 12'b111111111111;
assign CPM[9230] = 12'b111111111111;
assign CPM[9231] = 12'b111111111111;
assign CPM[9232] = 12'b111111111111;
assign CPM[9233] = 12'b111111111111;
assign CPM[9234] = 12'b111111111111;
assign CPM[9235] = 12'b111111111111;
assign CPM[9236] = 12'b111111111111;
assign CPM[9237] = 12'b111111111111;
assign CPM[9238] = 12'b111111111111;
assign CPM[9239] = 12'b111111111111;
assign CPM[9240] = 12'b111111111111;
assign CPM[9241] = 12'b111111111111;
assign CPM[9242] = 12'b111111111111;
assign CPM[9243] = 12'b111111111111;
assign CPM[9244] = 12'b111111111111;
assign CPM[9245] = 12'b111111111111;
assign CPM[9246] = 12'b111111111111;
assign CPM[9247] = 12'b111111111111;
assign CPM[9248] = 12'b111111111111;
assign CPM[9249] = 12'b111111111111;
assign CPM[9250] = 12'b111111111111;
assign CPM[9251] = 12'b111111111111;
assign CPM[9252] = 12'b111111111111;
assign CPM[9253] = 12'b111111111111;
assign CPM[9254] = 12'b111111111111;
assign CPM[9255] = 12'b111111111111;
assign CPM[9256] = 12'b111111111111;
assign CPM[9257] = 12'b111111111111;
assign CPM[9258] = 12'b111111111111;
assign CPM[9259] = 12'b111111111111;
assign CPM[9260] = 12'b111111111111;
assign CPM[9261] = 12'b111111111111;
assign CPM[9262] = 12'b111111111111;
assign CPM[9263] = 12'b111111111111;
assign CPM[9264] = 12'b111111111111;
assign CPM[9265] = 12'b111111111111;
assign CPM[9266] = 12'b111111111111;
assign CPM[9267] = 12'b111111111111;
assign CPM[9268] = 12'b111111111111;
assign CPM[9269] = 12'b111111111111;
assign CPM[9270] = 12'b111111111111;
assign CPM[9271] = 12'b111111111111;
assign CPM[9272] = 12'b111111111111;
assign CPM[9273] = 12'b111111111111;
assign CPM[9274] = 12'b111111111111;
assign CPM[9275] = 12'b111111111111;
assign CPM[9276] = 12'b111111111111;
assign CPM[9277] = 12'b111111111111;
assign CPM[9278] = 12'b111111111111;
assign CPM[9279] = 12'b111111111111;
assign CPM[9280] = 12'b111111111111;
assign CPM[9281] = 12'b111111111111;
assign CPM[9282] = 12'b111111111111;
assign CPM[9283] = 12'b111111111111;
assign CPM[9284] = 12'b111111111111;
assign CPM[9285] = 12'b111111111111;
assign CPM[9286] = 12'b111111111111;
assign CPM[9287] = 12'b111111111111;
assign CPM[9288] = 12'b111111111111;
assign CPM[9289] = 12'b111111111111;
assign CPM[9290] = 12'b111111111111;
assign CPM[9291] = 12'b111111111111;
assign CPM[9292] = 12'b111111111111;
assign CPM[9293] = 12'b111111111111;
assign CPM[9294] = 12'b111111111111;
assign CPM[9295] = 12'b111111111111;
assign CPM[9296] = 12'b111111111111;
assign CPM[9297] = 12'b111111111111;
assign CPM[9298] = 12'b111111111111;
assign CPM[9299] = 12'b111111111111;
assign CPM[9300] = 12'b111111111111;
assign CPM[9301] = 12'b111111111111;
assign CPM[9302] = 12'b111111111111;
assign CPM[9303] = 12'b111111111111;
assign CPM[9304] = 12'b111111111111;
assign CPM[9305] = 12'b111111111111;
assign CPM[9306] = 12'b111111111111;
assign CPM[9307] = 12'b111111111111;
assign CPM[9308] = 12'b111111111111;
assign CPM[9309] = 12'b111111111111;
assign CPM[9310] = 12'b111111111111;
assign CPM[9311] = 12'b111111111111;
assign CPM[9312] = 12'b111111111111;
assign CPM[9313] = 12'b111111111111;
assign CPM[9314] = 12'b111111111111;
assign CPM[9315] = 12'b111111111111;
assign CPM[9316] = 12'b111111111111;
assign CPM[9317] = 12'b111111111111;
assign CPM[9318] = 12'b111111111111;
assign CPM[9319] = 12'b111111111111;
assign CPM[9320] = 12'b111111111111;
assign CPM[9321] = 12'b000000000000;
assign CPM[9322] = 12'b000000000000;
assign CPM[9323] = 12'b000000000000;
assign CPM[9324] = 12'b000000000000;
assign CPM[9325] = 12'b000000000000;
assign CPM[9326] = 12'b000000000000;
assign CPM[9327] = 12'b000000000000;
assign CPM[9328] = 12'b000000000000;
assign CPM[9329] = 12'b000000000000;
assign CPM[9330] = 12'b000000000000;
assign CPM[9331] = 12'b000000000000;
assign CPM[9332] = 12'b000000000000;
assign CPM[9333] = 12'b000000000000;
assign CPM[9334] = 12'b000000000000;
assign CPM[9335] = 12'b111111111111;
assign CPM[9336] = 12'b111111111111;
assign CPM[9337] = 12'b111111111111;
assign CPM[9338] = 12'b111111111111;
assign CPM[9339] = 12'b111111111111;
assign CPM[9340] = 12'b111111111111;
assign CPM[9341] = 12'b111111111111;
assign CPM[9342] = 12'b111111111111;
assign CPM[9343] = 12'b111111111111;
assign CPM[9344] = 12'b111111111111;
assign CPM[9345] = 12'b111111111111;
assign CPM[9346] = 12'b111111111111;
assign CPM[9347] = 12'b111111111111;
assign CPM[9348] = 12'b111111111111;
assign CPM[9349] = 12'b111111111111;
assign CPM[9350] = 12'b111111111111;
assign CPM[9351] = 12'b111111111111;
assign CPM[9352] = 12'b111111111111;
assign CPM[9353] = 12'b000000000000;
assign CPM[9354] = 12'b000000000000;
assign CPM[9355] = 12'b000000000000;
assign CPM[9356] = 12'b000000000000;
assign CPM[9357] = 12'b000000000000;
assign CPM[9358] = 12'b000000000000;
assign CPM[9359] = 12'b000000000000;
assign CPM[9360] = 12'b000000000000;
assign CPM[9361] = 12'b000000000000;
assign CPM[9362] = 12'b000000000000;
assign CPM[9363] = 12'b000000000000;
assign CPM[9364] = 12'b000000000000;
assign CPM[9365] = 12'b000000000000;
assign CPM[9366] = 12'b000000000000;
assign CPM[9367] = 12'b111111111111;
assign CPM[9368] = 12'b111111111111;
assign CPM[9369] = 12'b111111111111;
assign CPM[9370] = 12'b111111111111;
assign CPM[9371] = 12'b111111111111;
assign CPM[9372] = 12'b111111111111;
assign CPM[9373] = 12'b111111111111;
assign CPM[9374] = 12'b111111111111;
assign CPM[9375] = 12'b111111111111;
assign CPM[9376] = 12'b111111111111;
assign CPM[9377] = 12'b111111111111;
assign CPM[9378] = 12'b111111111111;
assign CPM[9379] = 12'b111111111111;
assign CPM[9380] = 12'b111111111111;
assign CPM[9381] = 12'b111111111111;
assign CPM[9382] = 12'b111111111111;
assign CPM[9383] = 12'b111111111111;
assign CPM[9384] = 12'b111111111111;
assign CPM[9385] = 12'b000000000000;
assign CPM[9386] = 12'b000000000000;
assign CPM[9387] = 12'b000000000000;
assign CPM[9388] = 12'b000000000000;
assign CPM[9389] = 12'b000000000000;
assign CPM[9390] = 12'b000000000000;
assign CPM[9391] = 12'b000000000000;
assign CPM[9392] = 12'b000000000000;
assign CPM[9393] = 12'b000000000000;
assign CPM[9394] = 12'b000000000000;
assign CPM[9395] = 12'b000000000000;
assign CPM[9396] = 12'b000000000000;
assign CPM[9397] = 12'b000000000000;
assign CPM[9398] = 12'b000000000000;
assign CPM[9399] = 12'b111111111111;
assign CPM[9400] = 12'b111111111111;
assign CPM[9401] = 12'b111111111111;
assign CPM[9402] = 12'b111111111111;
assign CPM[9403] = 12'b111111111111;
assign CPM[9404] = 12'b111111111111;
assign CPM[9405] = 12'b111111111111;
assign CPM[9406] = 12'b111111111111;
assign CPM[9407] = 12'b111111111111;
assign CPM[9408] = 12'b111111111111;
assign CPM[9409] = 12'b111111111111;
assign CPM[9410] = 12'b111111111111;
assign CPM[9411] = 12'b111111111111;
assign CPM[9412] = 12'b111111111111;
assign CPM[9413] = 12'b111111111111;
assign CPM[9414] = 12'b111111111111;
assign CPM[9415] = 12'b111111111111;
assign CPM[9416] = 12'b111111111111;
assign CPM[9417] = 12'b000000000000;
assign CPM[9418] = 12'b000000000000;
assign CPM[9419] = 12'b000000000000;
assign CPM[9420] = 12'b000000000000;
assign CPM[9421] = 12'b000000000000;
assign CPM[9422] = 12'b000000000000;
assign CPM[9423] = 12'b000000000000;
assign CPM[9424] = 12'b000000000000;
assign CPM[9425] = 12'b000000000000;
assign CPM[9426] = 12'b000000000000;
assign CPM[9427] = 12'b000000000000;
assign CPM[9428] = 12'b000000000000;
assign CPM[9429] = 12'b000000000000;
assign CPM[9430] = 12'b000000000000;
assign CPM[9431] = 12'b111111111111;
assign CPM[9432] = 12'b111111111111;
assign CPM[9433] = 12'b111111111111;
assign CPM[9434] = 12'b111111111111;
assign CPM[9435] = 12'b111111111111;
assign CPM[9436] = 12'b111111111111;
assign CPM[9437] = 12'b111111111111;
assign CPM[9438] = 12'b111111111111;
assign CPM[9439] = 12'b111111111111;
assign CPM[9440] = 12'b111111111111;
assign CPM[9441] = 12'b111111111111;
assign CPM[9442] = 12'b111111111111;
assign CPM[9443] = 12'b111111111111;
assign CPM[9444] = 12'b111111111111;
assign CPM[9445] = 12'b000000000000;
assign CPM[9446] = 12'b000000000000;
assign CPM[9447] = 12'b000000000000;
assign CPM[9448] = 12'b000000000000;
assign CPM[9449] = 12'b111111111111;
assign CPM[9450] = 12'b111111111111;
assign CPM[9451] = 12'b111111111111;
assign CPM[9452] = 12'b111111111111;
assign CPM[9453] = 12'b111111111111;
assign CPM[9454] = 12'b111111111111;
assign CPM[9455] = 12'b111111111111;
assign CPM[9456] = 12'b111111111111;
assign CPM[9457] = 12'b111111111111;
assign CPM[9458] = 12'b111111111111;
assign CPM[9459] = 12'b111111111111;
assign CPM[9460] = 12'b111111111111;
assign CPM[9461] = 12'b111111111111;
assign CPM[9462] = 12'b111111111111;
assign CPM[9463] = 12'b111111111111;
assign CPM[9464] = 12'b111111111111;
assign CPM[9465] = 12'b111111111111;
assign CPM[9466] = 12'b111111111111;
assign CPM[9467] = 12'b111111111111;
assign CPM[9468] = 12'b111111111111;
assign CPM[9469] = 12'b111111111111;
assign CPM[9470] = 12'b111111111111;
assign CPM[9471] = 12'b111111111111;
assign CPM[9472] = 12'b111111111111;
assign CPM[9473] = 12'b111111111111;
assign CPM[9474] = 12'b111111111111;
assign CPM[9475] = 12'b111111111111;
assign CPM[9476] = 12'b111111111111;
assign CPM[9477] = 12'b000000000000;
assign CPM[9478] = 12'b000000000000;
assign CPM[9479] = 12'b000000000000;
assign CPM[9480] = 12'b000000000000;
assign CPM[9481] = 12'b111111111111;
assign CPM[9482] = 12'b111111111111;
assign CPM[9483] = 12'b111111111111;
assign CPM[9484] = 12'b111111111111;
assign CPM[9485] = 12'b111111111111;
assign CPM[9486] = 12'b111111111111;
assign CPM[9487] = 12'b111111111111;
assign CPM[9488] = 12'b111111111111;
assign CPM[9489] = 12'b111111111111;
assign CPM[9490] = 12'b111111111111;
assign CPM[9491] = 12'b111111111111;
assign CPM[9492] = 12'b111111111111;
assign CPM[9493] = 12'b111111111111;
assign CPM[9494] = 12'b111111111111;
assign CPM[9495] = 12'b111111111111;
assign CPM[9496] = 12'b111111111111;
assign CPM[9497] = 12'b111111111111;
assign CPM[9498] = 12'b111111111111;
assign CPM[9499] = 12'b111111111111;
assign CPM[9500] = 12'b111111111111;
assign CPM[9501] = 12'b111111111111;
assign CPM[9502] = 12'b111111111111;
assign CPM[9503] = 12'b111111111111;
assign CPM[9504] = 12'b111111111111;
assign CPM[9505] = 12'b111111111111;
assign CPM[9506] = 12'b111111111111;
assign CPM[9507] = 12'b111111111111;
assign CPM[9508] = 12'b111111111111;
assign CPM[9509] = 12'b000000000000;
assign CPM[9510] = 12'b000000000000;
assign CPM[9511] = 12'b000000000000;
assign CPM[9512] = 12'b000000000000;
assign CPM[9513] = 12'b111111111111;
assign CPM[9514] = 12'b111111111111;
assign CPM[9515] = 12'b111111111111;
assign CPM[9516] = 12'b111111111111;
assign CPM[9517] = 12'b111111111111;
assign CPM[9518] = 12'b111111111111;
assign CPM[9519] = 12'b111111111111;
assign CPM[9520] = 12'b111111111111;
assign CPM[9521] = 12'b111111111111;
assign CPM[9522] = 12'b111111111111;
assign CPM[9523] = 12'b111111111111;
assign CPM[9524] = 12'b111111111111;
assign CPM[9525] = 12'b111111111111;
assign CPM[9526] = 12'b111111111111;
assign CPM[9527] = 12'b111111111111;
assign CPM[9528] = 12'b111111111111;
assign CPM[9529] = 12'b111111111111;
assign CPM[9530] = 12'b111111111111;
assign CPM[9531] = 12'b111111111111;
assign CPM[9532] = 12'b111111111111;
assign CPM[9533] = 12'b111111111111;
assign CPM[9534] = 12'b111111111111;
assign CPM[9535] = 12'b111111111111;
assign CPM[9536] = 12'b111111111111;
assign CPM[9537] = 12'b111111111111;
assign CPM[9538] = 12'b111111111111;
assign CPM[9539] = 12'b111111111111;
assign CPM[9540] = 12'b111111111111;
assign CPM[9541] = 12'b000000000000;
assign CPM[9542] = 12'b000000000000;
assign CPM[9543] = 12'b000000000000;
assign CPM[9544] = 12'b000000000000;
assign CPM[9545] = 12'b111111111111;
assign CPM[9546] = 12'b111111111111;
assign CPM[9547] = 12'b111111111111;
assign CPM[9548] = 12'b111111111111;
assign CPM[9549] = 12'b111111111111;
assign CPM[9550] = 12'b111111111111;
assign CPM[9551] = 12'b111111111111;
assign CPM[9552] = 12'b111111111111;
assign CPM[9553] = 12'b111111111111;
assign CPM[9554] = 12'b111111111111;
assign CPM[9555] = 12'b111111111111;
assign CPM[9556] = 12'b111111111111;
assign CPM[9557] = 12'b111111111111;
assign CPM[9558] = 12'b111111111111;
assign CPM[9559] = 12'b111111111111;
assign CPM[9560] = 12'b111111111111;
assign CPM[9561] = 12'b111111111111;
assign CPM[9562] = 12'b111111111111;
assign CPM[9563] = 12'b111111111111;
assign CPM[9564] = 12'b111111111111;
assign CPM[9565] = 12'b111111111111;
assign CPM[9566] = 12'b111111111111;
assign CPM[9567] = 12'b111111111111;
assign CPM[9568] = 12'b111111111111;
assign CPM[9569] = 12'b111111111111;
assign CPM[9570] = 12'b111111111111;
assign CPM[9571] = 12'b111111111111;
assign CPM[9572] = 12'b111111111111;
assign CPM[9573] = 12'b000000000000;
assign CPM[9574] = 12'b000000000000;
assign CPM[9575] = 12'b000000000000;
assign CPM[9576] = 12'b000000000000;
assign CPM[9577] = 12'b111111111111;
assign CPM[9578] = 12'b111111111111;
assign CPM[9579] = 12'b111111111111;
assign CPM[9580] = 12'b111111111111;
assign CPM[9581] = 12'b111111111111;
assign CPM[9582] = 12'b111111111111;
assign CPM[9583] = 12'b111111111111;
assign CPM[9584] = 12'b111111111111;
assign CPM[9585] = 12'b111111111111;
assign CPM[9586] = 12'b111111111111;
assign CPM[9587] = 12'b111111111111;
assign CPM[9588] = 12'b111111111111;
assign CPM[9589] = 12'b111111111111;
assign CPM[9590] = 12'b111111111111;
assign CPM[9591] = 12'b111111111111;
assign CPM[9592] = 12'b111111111111;
assign CPM[9593] = 12'b111111111111;
assign CPM[9594] = 12'b111111111111;
assign CPM[9595] = 12'b111111111111;
assign CPM[9596] = 12'b111111111111;
assign CPM[9597] = 12'b111111111111;
assign CPM[9598] = 12'b111111111111;
assign CPM[9599] = 12'b111111111111;
assign CPM[9600] = 12'b111111111111;
assign CPM[9601] = 12'b111111111111;
assign CPM[9602] = 12'b111111111111;
assign CPM[9603] = 12'b111111111111;
assign CPM[9604] = 12'b111111111111;
assign CPM[9605] = 12'b000000000000;
assign CPM[9606] = 12'b000000000000;
assign CPM[9607] = 12'b000000000000;
assign CPM[9608] = 12'b000000000000;
assign CPM[9609] = 12'b111111111111;
assign CPM[9610] = 12'b111111111111;
assign CPM[9611] = 12'b111111111111;
assign CPM[9612] = 12'b111111111111;
assign CPM[9613] = 12'b111111111111;
assign CPM[9614] = 12'b111111111111;
assign CPM[9615] = 12'b111111111111;
assign CPM[9616] = 12'b111111111111;
assign CPM[9617] = 12'b111111111111;
assign CPM[9618] = 12'b111111111111;
assign CPM[9619] = 12'b111111111111;
assign CPM[9620] = 12'b111111111111;
assign CPM[9621] = 12'b111111111111;
assign CPM[9622] = 12'b111111111111;
assign CPM[9623] = 12'b111111111111;
assign CPM[9624] = 12'b111111111111;
assign CPM[9625] = 12'b111111111111;
assign CPM[9626] = 12'b111111111111;
assign CPM[9627] = 12'b111111111111;
assign CPM[9628] = 12'b111111111111;
assign CPM[9629] = 12'b111111111111;
assign CPM[9630] = 12'b111111111111;
assign CPM[9631] = 12'b111111111111;
assign CPM[9632] = 12'b111111111111;
assign CPM[9633] = 12'b111111111111;
assign CPM[9634] = 12'b111111111111;
assign CPM[9635] = 12'b111111111111;
assign CPM[9636] = 12'b111111111111;
assign CPM[9637] = 12'b000000000000;
assign CPM[9638] = 12'b000000000000;
assign CPM[9639] = 12'b000000000000;
assign CPM[9640] = 12'b000000000000;
assign CPM[9641] = 12'b111111111111;
assign CPM[9642] = 12'b111111111111;
assign CPM[9643] = 12'b111111111111;
assign CPM[9644] = 12'b111111111111;
assign CPM[9645] = 12'b111111111111;
assign CPM[9646] = 12'b111111111111;
assign CPM[9647] = 12'b111111111111;
assign CPM[9648] = 12'b111111111111;
assign CPM[9649] = 12'b111111111111;
assign CPM[9650] = 12'b111111111111;
assign CPM[9651] = 12'b111111111111;
assign CPM[9652] = 12'b111111111111;
assign CPM[9653] = 12'b111111111111;
assign CPM[9654] = 12'b111111111111;
assign CPM[9655] = 12'b111111111111;
assign CPM[9656] = 12'b111111111111;
assign CPM[9657] = 12'b111111111111;
assign CPM[9658] = 12'b111111111111;
assign CPM[9659] = 12'b111111111111;
assign CPM[9660] = 12'b111111111111;
assign CPM[9661] = 12'b111111111111;
assign CPM[9662] = 12'b111111111111;
assign CPM[9663] = 12'b111111111111;
assign CPM[9664] = 12'b111111111111;
assign CPM[9665] = 12'b111111111111;
assign CPM[9666] = 12'b111111111111;
assign CPM[9667] = 12'b111111111111;
assign CPM[9668] = 12'b111111111111;
assign CPM[9669] = 12'b000000000000;
assign CPM[9670] = 12'b000000000000;
assign CPM[9671] = 12'b000000000000;
assign CPM[9672] = 12'b000000000000;
assign CPM[9673] = 12'b000000000000;
assign CPM[9674] = 12'b000000000000;
assign CPM[9675] = 12'b000000000000;
assign CPM[9676] = 12'b000000000000;
assign CPM[9677] = 12'b000000000000;
assign CPM[9678] = 12'b000000000000;
assign CPM[9679] = 12'b000000000000;
assign CPM[9680] = 12'b000000000000;
assign CPM[9681] = 12'b000000000000;
assign CPM[9682] = 12'b000000000000;
assign CPM[9683] = 12'b000000000000;
assign CPM[9684] = 12'b000000000000;
assign CPM[9685] = 12'b111111111111;
assign CPM[9686] = 12'b111111111111;
assign CPM[9687] = 12'b111111111111;
assign CPM[9688] = 12'b111111111111;
assign CPM[9689] = 12'b111111111111;
assign CPM[9690] = 12'b111111111111;
assign CPM[9691] = 12'b111111111111;
assign CPM[9692] = 12'b111111111111;
assign CPM[9693] = 12'b111111111111;
assign CPM[9694] = 12'b111111111111;
assign CPM[9695] = 12'b111111111111;
assign CPM[9696] = 12'b111111111111;
assign CPM[9697] = 12'b111111111111;
assign CPM[9698] = 12'b111111111111;
assign CPM[9699] = 12'b111111111111;
assign CPM[9700] = 12'b111111111111;
assign CPM[9701] = 12'b000000000000;
assign CPM[9702] = 12'b000000000000;
assign CPM[9703] = 12'b000000000000;
assign CPM[9704] = 12'b000000000000;
assign CPM[9705] = 12'b000000000000;
assign CPM[9706] = 12'b000000000000;
assign CPM[9707] = 12'b000000000000;
assign CPM[9708] = 12'b000000000000;
assign CPM[9709] = 12'b000000000000;
assign CPM[9710] = 12'b000000000000;
assign CPM[9711] = 12'b000000000000;
assign CPM[9712] = 12'b000000000000;
assign CPM[9713] = 12'b000000000000;
assign CPM[9714] = 12'b000000000000;
assign CPM[9715] = 12'b000000000000;
assign CPM[9716] = 12'b000000000000;
assign CPM[9717] = 12'b111111111111;
assign CPM[9718] = 12'b111111111111;
assign CPM[9719] = 12'b111111111111;
assign CPM[9720] = 12'b111111111111;
assign CPM[9721] = 12'b111111111111;
assign CPM[9722] = 12'b111111111111;
assign CPM[9723] = 12'b111111111111;
assign CPM[9724] = 12'b111111111111;
assign CPM[9725] = 12'b111111111111;
assign CPM[9726] = 12'b111111111111;
assign CPM[9727] = 12'b111111111111;
assign CPM[9728] = 12'b111111111111;
assign CPM[9729] = 12'b111111111111;
assign CPM[9730] = 12'b111111111111;
assign CPM[9731] = 12'b111111111111;
assign CPM[9732] = 12'b111111111111;
assign CPM[9733] = 12'b000000000000;
assign CPM[9734] = 12'b000000000000;
assign CPM[9735] = 12'b000000000000;
assign CPM[9736] = 12'b000000000000;
assign CPM[9737] = 12'b000000000000;
assign CPM[9738] = 12'b000000000000;
assign CPM[9739] = 12'b000000000000;
assign CPM[9740] = 12'b000000000000;
assign CPM[9741] = 12'b000000000000;
assign CPM[9742] = 12'b000000000000;
assign CPM[9743] = 12'b000000000000;
assign CPM[9744] = 12'b000000000000;
assign CPM[9745] = 12'b000000000000;
assign CPM[9746] = 12'b000000000000;
assign CPM[9747] = 12'b000000000000;
assign CPM[9748] = 12'b000000000000;
assign CPM[9749] = 12'b111111111111;
assign CPM[9750] = 12'b111111111111;
assign CPM[9751] = 12'b111111111111;
assign CPM[9752] = 12'b111111111111;
assign CPM[9753] = 12'b111111111111;
assign CPM[9754] = 12'b111111111111;
assign CPM[9755] = 12'b111111111111;
assign CPM[9756] = 12'b111111111111;
assign CPM[9757] = 12'b111111111111;
assign CPM[9758] = 12'b111111111111;
assign CPM[9759] = 12'b111111111111;
assign CPM[9760] = 12'b111111111111;
assign CPM[9761] = 12'b111111111111;
assign CPM[9762] = 12'b111111111111;
assign CPM[9763] = 12'b111111111111;
assign CPM[9764] = 12'b111111111111;
assign CPM[9765] = 12'b000000000000;
assign CPM[9766] = 12'b000000000000;
assign CPM[9767] = 12'b000000000000;
assign CPM[9768] = 12'b000000000000;
assign CPM[9769] = 12'b000000000000;
assign CPM[9770] = 12'b000000000000;
assign CPM[9771] = 12'b000000000000;
assign CPM[9772] = 12'b000000000000;
assign CPM[9773] = 12'b000000000000;
assign CPM[9774] = 12'b000000000000;
assign CPM[9775] = 12'b000000000000;
assign CPM[9776] = 12'b000000000000;
assign CPM[9777] = 12'b000000000000;
assign CPM[9778] = 12'b000000000000;
assign CPM[9779] = 12'b000000000000;
assign CPM[9780] = 12'b000000000000;
assign CPM[9781] = 12'b111111111111;
assign CPM[9782] = 12'b111111111111;
assign CPM[9783] = 12'b111111111111;
assign CPM[9784] = 12'b111111111111;
assign CPM[9785] = 12'b111111111111;
assign CPM[9786] = 12'b111111111111;
assign CPM[9787] = 12'b111111111111;
assign CPM[9788] = 12'b111111111111;
assign CPM[9789] = 12'b111111111111;
assign CPM[9790] = 12'b111111111111;
assign CPM[9791] = 12'b111111111111;
assign CPM[9792] = 12'b111111111111;
assign CPM[9793] = 12'b111111111111;
assign CPM[9794] = 12'b111111111111;
assign CPM[9795] = 12'b111111111111;
assign CPM[9796] = 12'b111111111111;
assign CPM[9797] = 12'b000000000000;
assign CPM[9798] = 12'b000000000000;
assign CPM[9799] = 12'b000000000000;
assign CPM[9800] = 12'b000000000000;
assign CPM[9801] = 12'b111111111111;
assign CPM[9802] = 12'b111111111111;
assign CPM[9803] = 12'b111111111111;
assign CPM[9804] = 12'b111111111111;
assign CPM[9805] = 12'b111111111111;
assign CPM[9806] = 12'b111111111111;
assign CPM[9807] = 12'b111111111111;
assign CPM[9808] = 12'b111111111111;
assign CPM[9809] = 12'b111111111111;
assign CPM[9810] = 12'b111111111111;
assign CPM[9811] = 12'b111111111111;
assign CPM[9812] = 12'b111111111111;
assign CPM[9813] = 12'b000000000000;
assign CPM[9814] = 12'b000000000000;
assign CPM[9815] = 12'b000000000000;
assign CPM[9816] = 12'b000000000000;
assign CPM[9817] = 12'b111111111111;
assign CPM[9818] = 12'b111111111111;
assign CPM[9819] = 12'b111111111111;
assign CPM[9820] = 12'b111111111111;
assign CPM[9821] = 12'b111111111111;
assign CPM[9822] = 12'b111111111111;
assign CPM[9823] = 12'b111111111111;
assign CPM[9824] = 12'b111111111111;
assign CPM[9825] = 12'b111111111111;
assign CPM[9826] = 12'b111111111111;
assign CPM[9827] = 12'b111111111111;
assign CPM[9828] = 12'b111111111111;
assign CPM[9829] = 12'b000000000000;
assign CPM[9830] = 12'b000000000000;
assign CPM[9831] = 12'b000000000000;
assign CPM[9832] = 12'b000000000000;
assign CPM[9833] = 12'b111111111111;
assign CPM[9834] = 12'b111111111111;
assign CPM[9835] = 12'b111111111111;
assign CPM[9836] = 12'b111111111111;
assign CPM[9837] = 12'b111111111111;
assign CPM[9838] = 12'b111111111111;
assign CPM[9839] = 12'b111111111111;
assign CPM[9840] = 12'b111111111111;
assign CPM[9841] = 12'b111111111111;
assign CPM[9842] = 12'b111111111111;
assign CPM[9843] = 12'b111111111111;
assign CPM[9844] = 12'b111111111111;
assign CPM[9845] = 12'b000000000000;
assign CPM[9846] = 12'b000000000000;
assign CPM[9847] = 12'b000000000000;
assign CPM[9848] = 12'b000000000000;
assign CPM[9849] = 12'b111111111111;
assign CPM[9850] = 12'b111111111111;
assign CPM[9851] = 12'b111111111111;
assign CPM[9852] = 12'b111111111111;
assign CPM[9853] = 12'b111111111111;
assign CPM[9854] = 12'b111111111111;
assign CPM[9855] = 12'b111111111111;
assign CPM[9856] = 12'b111111111111;
assign CPM[9857] = 12'b111111111111;
assign CPM[9858] = 12'b111111111111;
assign CPM[9859] = 12'b111111111111;
assign CPM[9860] = 12'b111111111111;
assign CPM[9861] = 12'b000000000000;
assign CPM[9862] = 12'b000000000000;
assign CPM[9863] = 12'b000000000000;
assign CPM[9864] = 12'b000000000000;
assign CPM[9865] = 12'b111111111111;
assign CPM[9866] = 12'b111111111111;
assign CPM[9867] = 12'b111111111111;
assign CPM[9868] = 12'b111111111111;
assign CPM[9869] = 12'b111111111111;
assign CPM[9870] = 12'b111111111111;
assign CPM[9871] = 12'b111111111111;
assign CPM[9872] = 12'b111111111111;
assign CPM[9873] = 12'b111111111111;
assign CPM[9874] = 12'b111111111111;
assign CPM[9875] = 12'b111111111111;
assign CPM[9876] = 12'b111111111111;
assign CPM[9877] = 12'b000000000000;
assign CPM[9878] = 12'b000000000000;
assign CPM[9879] = 12'b000000000000;
assign CPM[9880] = 12'b000000000000;
assign CPM[9881] = 12'b111111111111;
assign CPM[9882] = 12'b111111111111;
assign CPM[9883] = 12'b111111111111;
assign CPM[9884] = 12'b111111111111;
assign CPM[9885] = 12'b111111111111;
assign CPM[9886] = 12'b111111111111;
assign CPM[9887] = 12'b111111111111;
assign CPM[9888] = 12'b111111111111;
assign CPM[9889] = 12'b111111111111;
assign CPM[9890] = 12'b111111111111;
assign CPM[9891] = 12'b111111111111;
assign CPM[9892] = 12'b111111111111;
assign CPM[9893] = 12'b000000000000;
assign CPM[9894] = 12'b000000000000;
assign CPM[9895] = 12'b000000000000;
assign CPM[9896] = 12'b000000000000;
assign CPM[9897] = 12'b111111111111;
assign CPM[9898] = 12'b111111111111;
assign CPM[9899] = 12'b111111111111;
assign CPM[9900] = 12'b111111111111;
assign CPM[9901] = 12'b111111111111;
assign CPM[9902] = 12'b111111111111;
assign CPM[9903] = 12'b111111111111;
assign CPM[9904] = 12'b111111111111;
assign CPM[9905] = 12'b111111111111;
assign CPM[9906] = 12'b111111111111;
assign CPM[9907] = 12'b111111111111;
assign CPM[9908] = 12'b111111111111;
assign CPM[9909] = 12'b000000000000;
assign CPM[9910] = 12'b000000000000;
assign CPM[9911] = 12'b000000000000;
assign CPM[9912] = 12'b000000000000;
assign CPM[9913] = 12'b111111111111;
assign CPM[9914] = 12'b111111111111;
assign CPM[9915] = 12'b111111111111;
assign CPM[9916] = 12'b111111111111;
assign CPM[9917] = 12'b111111111111;
assign CPM[9918] = 12'b111111111111;
assign CPM[9919] = 12'b111111111111;
assign CPM[9920] = 12'b111111111111;
assign CPM[9921] = 12'b111111111111;
assign CPM[9922] = 12'b111111111111;
assign CPM[9923] = 12'b111111111111;
assign CPM[9924] = 12'b111111111111;
assign CPM[9925] = 12'b000000000000;
assign CPM[9926] = 12'b000000000000;
assign CPM[9927] = 12'b000000000000;
assign CPM[9928] = 12'b000000000000;
assign CPM[9929] = 12'b111111111111;
assign CPM[9930] = 12'b111111111111;
assign CPM[9931] = 12'b111111111111;
assign CPM[9932] = 12'b111111111111;
assign CPM[9933] = 12'b111111111111;
assign CPM[9934] = 12'b111111111111;
assign CPM[9935] = 12'b111111111111;
assign CPM[9936] = 12'b111111111111;
assign CPM[9937] = 12'b111111111111;
assign CPM[9938] = 12'b111111111111;
assign CPM[9939] = 12'b111111111111;
assign CPM[9940] = 12'b111111111111;
assign CPM[9941] = 12'b000000000000;
assign CPM[9942] = 12'b000000000000;
assign CPM[9943] = 12'b000000000000;
assign CPM[9944] = 12'b000000000000;
assign CPM[9945] = 12'b111111111111;
assign CPM[9946] = 12'b111111111111;
assign CPM[9947] = 12'b111111111111;
assign CPM[9948] = 12'b111111111111;
assign CPM[9949] = 12'b111111111111;
assign CPM[9950] = 12'b111111111111;
assign CPM[9951] = 12'b111111111111;
assign CPM[9952] = 12'b111111111111;
assign CPM[9953] = 12'b111111111111;
assign CPM[9954] = 12'b111111111111;
assign CPM[9955] = 12'b111111111111;
assign CPM[9956] = 12'b111111111111;
assign CPM[9957] = 12'b000000000000;
assign CPM[9958] = 12'b000000000000;
assign CPM[9959] = 12'b000000000000;
assign CPM[9960] = 12'b000000000000;
assign CPM[9961] = 12'b111111111111;
assign CPM[9962] = 12'b111111111111;
assign CPM[9963] = 12'b111111111111;
assign CPM[9964] = 12'b111111111111;
assign CPM[9965] = 12'b111111111111;
assign CPM[9966] = 12'b111111111111;
assign CPM[9967] = 12'b111111111111;
assign CPM[9968] = 12'b111111111111;
assign CPM[9969] = 12'b111111111111;
assign CPM[9970] = 12'b111111111111;
assign CPM[9971] = 12'b111111111111;
assign CPM[9972] = 12'b111111111111;
assign CPM[9973] = 12'b000000000000;
assign CPM[9974] = 12'b000000000000;
assign CPM[9975] = 12'b000000000000;
assign CPM[9976] = 12'b000000000000;
assign CPM[9977] = 12'b111111111111;
assign CPM[9978] = 12'b111111111111;
assign CPM[9979] = 12'b111111111111;
assign CPM[9980] = 12'b111111111111;
assign CPM[9981] = 12'b111111111111;
assign CPM[9982] = 12'b111111111111;
assign CPM[9983] = 12'b111111111111;
assign CPM[9984] = 12'b111111111111;
assign CPM[9985] = 12'b111111111111;
assign CPM[9986] = 12'b111111111111;
assign CPM[9987] = 12'b111111111111;
assign CPM[9988] = 12'b111111111111;
assign CPM[9989] = 12'b000000000000;
assign CPM[9990] = 12'b000000000000;
assign CPM[9991] = 12'b000000000000;
assign CPM[9992] = 12'b000000000000;
assign CPM[9993] = 12'b111111111111;
assign CPM[9994] = 12'b111111111111;
assign CPM[9995] = 12'b111111111111;
assign CPM[9996] = 12'b111111111111;
assign CPM[9997] = 12'b111111111111;
assign CPM[9998] = 12'b111111111111;
assign CPM[9999] = 12'b111111111111;
assign CPM[10000] = 12'b111111111111;
assign CPM[10001] = 12'b111111111111;
assign CPM[10002] = 12'b111111111111;
assign CPM[10003] = 12'b111111111111;
assign CPM[10004] = 12'b111111111111;
assign CPM[10005] = 12'b000000000000;
assign CPM[10006] = 12'b000000000000;
assign CPM[10007] = 12'b000000000000;
assign CPM[10008] = 12'b000000000000;
assign CPM[10009] = 12'b111111111111;
assign CPM[10010] = 12'b111111111111;
assign CPM[10011] = 12'b111111111111;
assign CPM[10012] = 12'b111111111111;
assign CPM[10013] = 12'b111111111111;
assign CPM[10014] = 12'b111111111111;
assign CPM[10015] = 12'b111111111111;
assign CPM[10016] = 12'b111111111111;
assign CPM[10017] = 12'b111111111111;
assign CPM[10018] = 12'b111111111111;
assign CPM[10019] = 12'b111111111111;
assign CPM[10020] = 12'b111111111111;
assign CPM[10021] = 12'b000000000000;
assign CPM[10022] = 12'b000000000000;
assign CPM[10023] = 12'b000000000000;
assign CPM[10024] = 12'b000000000000;
assign CPM[10025] = 12'b111111111111;
assign CPM[10026] = 12'b111111111111;
assign CPM[10027] = 12'b111111111111;
assign CPM[10028] = 12'b111111111111;
assign CPM[10029] = 12'b111111111111;
assign CPM[10030] = 12'b111111111111;
assign CPM[10031] = 12'b111111111111;
assign CPM[10032] = 12'b111111111111;
assign CPM[10033] = 12'b111111111111;
assign CPM[10034] = 12'b111111111111;
assign CPM[10035] = 12'b111111111111;
assign CPM[10036] = 12'b111111111111;
assign CPM[10037] = 12'b000000000000;
assign CPM[10038] = 12'b000000000000;
assign CPM[10039] = 12'b000000000000;
assign CPM[10040] = 12'b000000000000;
assign CPM[10041] = 12'b111111111111;
assign CPM[10042] = 12'b111111111111;
assign CPM[10043] = 12'b111111111111;
assign CPM[10044] = 12'b111111111111;
assign CPM[10045] = 12'b111111111111;
assign CPM[10046] = 12'b111111111111;
assign CPM[10047] = 12'b111111111111;
assign CPM[10048] = 12'b111111111111;
assign CPM[10049] = 12'b111111111111;
assign CPM[10050] = 12'b111111111111;
assign CPM[10051] = 12'b111111111111;
assign CPM[10052] = 12'b111111111111;
assign CPM[10053] = 12'b111111111111;
assign CPM[10054] = 12'b111111111111;
assign CPM[10055] = 12'b111111111111;
assign CPM[10056] = 12'b111111111111;
assign CPM[10057] = 12'b000000000000;
assign CPM[10058] = 12'b000000000000;
assign CPM[10059] = 12'b000000000000;
assign CPM[10060] = 12'b000000000000;
assign CPM[10061] = 12'b000000000000;
assign CPM[10062] = 12'b000000000000;
assign CPM[10063] = 12'b000000000000;
assign CPM[10064] = 12'b000000000000;
assign CPM[10065] = 12'b000000000000;
assign CPM[10066] = 12'b000000000000;
assign CPM[10067] = 12'b000000000000;
assign CPM[10068] = 12'b000000000000;
assign CPM[10069] = 12'b111111111111;
assign CPM[10070] = 12'b111111111111;
assign CPM[10071] = 12'b111111111111;
assign CPM[10072] = 12'b111111111111;
assign CPM[10073] = 12'b111111111111;
assign CPM[10074] = 12'b111111111111;
assign CPM[10075] = 12'b111111111111;
assign CPM[10076] = 12'b111111111111;
assign CPM[10077] = 12'b111111111111;
assign CPM[10078] = 12'b111111111111;
assign CPM[10079] = 12'b111111111111;
assign CPM[10080] = 12'b111111111111;
assign CPM[10081] = 12'b111111111111;
assign CPM[10082] = 12'b111111111111;
assign CPM[10083] = 12'b111111111111;
assign CPM[10084] = 12'b111111111111;
assign CPM[10085] = 12'b111111111111;
assign CPM[10086] = 12'b111111111111;
assign CPM[10087] = 12'b111111111111;
assign CPM[10088] = 12'b111111111111;
assign CPM[10089] = 12'b000000000000;
assign CPM[10090] = 12'b000000000000;
assign CPM[10091] = 12'b000000000000;
assign CPM[10092] = 12'b000000000000;
assign CPM[10093] = 12'b000000000000;
assign CPM[10094] = 12'b000000000000;
assign CPM[10095] = 12'b000000000000;
assign CPM[10096] = 12'b000000000000;
assign CPM[10097] = 12'b000000000000;
assign CPM[10098] = 12'b000000000000;
assign CPM[10099] = 12'b000000000000;
assign CPM[10100] = 12'b000000000000;
assign CPM[10101] = 12'b111111111111;
assign CPM[10102] = 12'b111111111111;
assign CPM[10103] = 12'b111111111111;
assign CPM[10104] = 12'b111111111111;
assign CPM[10105] = 12'b111111111111;
assign CPM[10106] = 12'b111111111111;
assign CPM[10107] = 12'b111111111111;
assign CPM[10108] = 12'b111111111111;
assign CPM[10109] = 12'b111111111111;
assign CPM[10110] = 12'b111111111111;
assign CPM[10111] = 12'b111111111111;
assign CPM[10112] = 12'b111111111111;
assign CPM[10113] = 12'b111111111111;
assign CPM[10114] = 12'b111111111111;
assign CPM[10115] = 12'b111111111111;
assign CPM[10116] = 12'b111111111111;
assign CPM[10117] = 12'b111111111111;
assign CPM[10118] = 12'b111111111111;
assign CPM[10119] = 12'b111111111111;
assign CPM[10120] = 12'b111111111111;
assign CPM[10121] = 12'b000000000000;
assign CPM[10122] = 12'b000000000000;
assign CPM[10123] = 12'b000000000000;
assign CPM[10124] = 12'b000000000000;
assign CPM[10125] = 12'b000000000000;
assign CPM[10126] = 12'b000000000000;
assign CPM[10127] = 12'b000000000000;
assign CPM[10128] = 12'b000000000000;
assign CPM[10129] = 12'b000000000000;
assign CPM[10130] = 12'b000000000000;
assign CPM[10131] = 12'b000000000000;
assign CPM[10132] = 12'b000000000000;
assign CPM[10133] = 12'b111111111111;
assign CPM[10134] = 12'b111111111111;
assign CPM[10135] = 12'b111111111111;
assign CPM[10136] = 12'b111111111111;
assign CPM[10137] = 12'b111111111111;
assign CPM[10138] = 12'b111111111111;
assign CPM[10139] = 12'b111111111111;
assign CPM[10140] = 12'b111111111111;
assign CPM[10141] = 12'b111111111111;
assign CPM[10142] = 12'b111111111111;
assign CPM[10143] = 12'b111111111111;
assign CPM[10144] = 12'b111111111111;
assign CPM[10145] = 12'b111111111111;
assign CPM[10146] = 12'b111111111111;
assign CPM[10147] = 12'b111111111111;
assign CPM[10148] = 12'b111111111111;
assign CPM[10149] = 12'b111111111111;
assign CPM[10150] = 12'b111111111111;
assign CPM[10151] = 12'b111111111111;
assign CPM[10152] = 12'b111111111111;
assign CPM[10153] = 12'b000000000000;
assign CPM[10154] = 12'b000000000000;
assign CPM[10155] = 12'b000000000000;
assign CPM[10156] = 12'b000000000000;
assign CPM[10157] = 12'b000000000000;
assign CPM[10158] = 12'b000000000000;
assign CPM[10159] = 12'b000000000000;
assign CPM[10160] = 12'b000000000000;
assign CPM[10161] = 12'b000000000000;
assign CPM[10162] = 12'b000000000000;
assign CPM[10163] = 12'b000000000000;
assign CPM[10164] = 12'b000000000000;
assign CPM[10165] = 12'b111111111111;
assign CPM[10166] = 12'b111111111111;
assign CPM[10167] = 12'b111111111111;
assign CPM[10168] = 12'b111111111111;
assign CPM[10169] = 12'b111111111111;
assign CPM[10170] = 12'b111111111111;
assign CPM[10171] = 12'b111111111111;
assign CPM[10172] = 12'b111111111111;
assign CPM[10173] = 12'b111111111111;
assign CPM[10174] = 12'b111111111111;
assign CPM[10175] = 12'b111111111111;
assign CPM[10176] = 12'b111111111111;
assign CPM[10177] = 12'b111111111111;
assign CPM[10178] = 12'b111111111111;
assign CPM[10179] = 12'b111111111111;
assign CPM[10180] = 12'b111111111111;
assign CPM[10181] = 12'b111111111111;
assign CPM[10182] = 12'b111111111111;
assign CPM[10183] = 12'b111111111111;
assign CPM[10184] = 12'b111111111111;
assign CPM[10185] = 12'b111111111111;
assign CPM[10186] = 12'b111111111111;
assign CPM[10187] = 12'b111111111111;
assign CPM[10188] = 12'b111111111111;
assign CPM[10189] = 12'b111111111111;
assign CPM[10190] = 12'b111111111111;
assign CPM[10191] = 12'b111111111111;
assign CPM[10192] = 12'b111111111111;
assign CPM[10193] = 12'b111111111111;
assign CPM[10194] = 12'b111111111111;
assign CPM[10195] = 12'b111111111111;
assign CPM[10196] = 12'b111111111111;
assign CPM[10197] = 12'b111111111111;
assign CPM[10198] = 12'b111111111111;
assign CPM[10199] = 12'b111111111111;
assign CPM[10200] = 12'b111111111111;
assign CPM[10201] = 12'b111111111111;
assign CPM[10202] = 12'b111111111111;
assign CPM[10203] = 12'b111111111111;
assign CPM[10204] = 12'b111111111111;
assign CPM[10205] = 12'b111111111111;
assign CPM[10206] = 12'b111111111111;
assign CPM[10207] = 12'b111111111111;
assign CPM[10208] = 12'b111111111111;
assign CPM[10209] = 12'b111111111111;
assign CPM[10210] = 12'b111111111111;
assign CPM[10211] = 12'b111111111111;
assign CPM[10212] = 12'b111111111111;
assign CPM[10213] = 12'b111111111111;
assign CPM[10214] = 12'b111111111111;
assign CPM[10215] = 12'b111111111111;
assign CPM[10216] = 12'b111111111111;
assign CPM[10217] = 12'b111111111111;
assign CPM[10218] = 12'b111111111111;
assign CPM[10219] = 12'b111111111111;
assign CPM[10220] = 12'b111111111111;
assign CPM[10221] = 12'b111111111111;
assign CPM[10222] = 12'b111111111111;
assign CPM[10223] = 12'b111111111111;
assign CPM[10224] = 12'b111111111111;
assign CPM[10225] = 12'b111111111111;
assign CPM[10226] = 12'b111111111111;
assign CPM[10227] = 12'b111111111111;
assign CPM[10228] = 12'b111111111111;
assign CPM[10229] = 12'b111111111111;
assign CPM[10230] = 12'b111111111111;
assign CPM[10231] = 12'b111111111111;
assign CPM[10232] = 12'b111111111111;
assign CPM[10233] = 12'b111111111111;
assign CPM[10234] = 12'b111111111111;
assign CPM[10235] = 12'b111111111111;
assign CPM[10236] = 12'b111111111111;
assign CPM[10237] = 12'b111111111111;
assign CPM[10238] = 12'b111111111111;
assign CPM[10239] = 12'b111111111111;
assign CPM[10240] = 12'b111111111111;
assign CPM[10241] = 12'b111111111111;
assign CPM[10242] = 12'b111111111111;
assign CPM[10243] = 12'b111111111111;
assign CPM[10244] = 12'b111111111111;
assign CPM[10245] = 12'b111111111111;
assign CPM[10246] = 12'b111111111111;
assign CPM[10247] = 12'b111111111111;
assign CPM[10248] = 12'b111111111111;
assign CPM[10249] = 12'b111111111111;
assign CPM[10250] = 12'b111111111111;
assign CPM[10251] = 12'b111111111111;
assign CPM[10252] = 12'b111111111111;
assign CPM[10253] = 12'b111111111111;
assign CPM[10254] = 12'b111111111111;
assign CPM[10255] = 12'b111111111111;
assign CPM[10256] = 12'b111111111111;
assign CPM[10257] = 12'b111111111111;
assign CPM[10258] = 12'b111111111111;
assign CPM[10259] = 12'b111111111111;
assign CPM[10260] = 12'b111111111111;
assign CPM[10261] = 12'b111111111111;
assign CPM[10262] = 12'b111111111111;
assign CPM[10263] = 12'b111111111111;
assign CPM[10264] = 12'b111111111111;
assign CPM[10265] = 12'b111111111111;
assign CPM[10266] = 12'b111111111111;
assign CPM[10267] = 12'b111111111111;
assign CPM[10268] = 12'b111111111111;
assign CPM[10269] = 12'b111111111111;
assign CPM[10270] = 12'b111111111111;
assign CPM[10271] = 12'b111111111111;
assign CPM[10272] = 12'b111111111111;
assign CPM[10273] = 12'b111111111111;
assign CPM[10274] = 12'b111111111111;
assign CPM[10275] = 12'b111111111111;
assign CPM[10276] = 12'b111111111111;
assign CPM[10277] = 12'b111111111111;
assign CPM[10278] = 12'b111111111111;
assign CPM[10279] = 12'b111111111111;
assign CPM[10280] = 12'b111111111111;
assign CPM[10281] = 12'b111111111111;
assign CPM[10282] = 12'b111111111111;
assign CPM[10283] = 12'b111111111111;
assign CPM[10284] = 12'b111111111111;
assign CPM[10285] = 12'b111111111111;
assign CPM[10286] = 12'b111111111111;
assign CPM[10287] = 12'b111111111111;
assign CPM[10288] = 12'b111111111111;
assign CPM[10289] = 12'b111111111111;
assign CPM[10290] = 12'b111111111111;
assign CPM[10291] = 12'b111111111111;
assign CPM[10292] = 12'b111111111111;
assign CPM[10293] = 12'b111111111111;
assign CPM[10294] = 12'b111111111111;
assign CPM[10295] = 12'b111111111111;
assign CPM[10296] = 12'b111111111111;
assign CPM[10297] = 12'b111111111111;
assign CPM[10298] = 12'b111111111111;
assign CPM[10299] = 12'b111111111111;
assign CPM[10300] = 12'b111111111111;
assign CPM[10301] = 12'b111111111111;
assign CPM[10302] = 12'b111111111111;
assign CPM[10303] = 12'b111111111111;
assign CPM[10304] = 12'b111111111111;
assign CPM[10305] = 12'b111111111111;
assign CPM[10306] = 12'b111111111111;
assign CPM[10307] = 12'b111111111111;
assign CPM[10308] = 12'b111111111111;
assign CPM[10309] = 12'b111111111111;
assign CPM[10310] = 12'b111111111111;
assign CPM[10311] = 12'b000000000000;
assign CPM[10312] = 12'b000000000000;
assign CPM[10313] = 12'b000000000000;
assign CPM[10314] = 12'b000000000000;
assign CPM[10315] = 12'b000000000000;
assign CPM[10316] = 12'b000000000000;
assign CPM[10317] = 12'b000000000000;
assign CPM[10318] = 12'b000000000000;
assign CPM[10319] = 12'b000000000000;
assign CPM[10320] = 12'b000000000000;
assign CPM[10321] = 12'b000000000000;
assign CPM[10322] = 12'b000000000000;
assign CPM[10323] = 12'b000000000000;
assign CPM[10324] = 12'b000000000000;
assign CPM[10325] = 12'b000000000000;
assign CPM[10326] = 12'b000000000000;
assign CPM[10327] = 12'b000000000000;
assign CPM[10328] = 12'b000000000000;
assign CPM[10329] = 12'b000000000000;
assign CPM[10330] = 12'b000000000000;
assign CPM[10331] = 12'b111111111111;
assign CPM[10332] = 12'b111111111111;
assign CPM[10333] = 12'b111111111111;
assign CPM[10334] = 12'b111111111111;
assign CPM[10335] = 12'b111111111111;
assign CPM[10336] = 12'b111111111111;
assign CPM[10337] = 12'b111111111111;
assign CPM[10338] = 12'b111111111111;
assign CPM[10339] = 12'b111111111111;
assign CPM[10340] = 12'b111111111111;
assign CPM[10341] = 12'b111111111111;
assign CPM[10342] = 12'b111111111111;
assign CPM[10343] = 12'b000000000000;
assign CPM[10344] = 12'b000000000000;
assign CPM[10345] = 12'b000000000000;
assign CPM[10346] = 12'b000000000000;
assign CPM[10347] = 12'b000000000000;
assign CPM[10348] = 12'b000000000000;
assign CPM[10349] = 12'b000000000000;
assign CPM[10350] = 12'b000000000000;
assign CPM[10351] = 12'b000000000000;
assign CPM[10352] = 12'b000000000000;
assign CPM[10353] = 12'b000000000000;
assign CPM[10354] = 12'b000000000000;
assign CPM[10355] = 12'b000000000000;
assign CPM[10356] = 12'b000000000000;
assign CPM[10357] = 12'b000000000000;
assign CPM[10358] = 12'b000000000000;
assign CPM[10359] = 12'b000000000000;
assign CPM[10360] = 12'b000000000000;
assign CPM[10361] = 12'b000000000000;
assign CPM[10362] = 12'b000000000000;
assign CPM[10363] = 12'b111111111111;
assign CPM[10364] = 12'b111111111111;
assign CPM[10365] = 12'b111111111111;
assign CPM[10366] = 12'b111111111111;
assign CPM[10367] = 12'b111111111111;
assign CPM[10368] = 12'b111111111111;
assign CPM[10369] = 12'b111111111111;
assign CPM[10370] = 12'b111111111111;
assign CPM[10371] = 12'b111111111111;
assign CPM[10372] = 12'b111111111111;
assign CPM[10373] = 12'b111111111111;
assign CPM[10374] = 12'b111111111111;
assign CPM[10375] = 12'b000000000000;
assign CPM[10376] = 12'b000000000000;
assign CPM[10377] = 12'b000000000000;
assign CPM[10378] = 12'b000000000000;
assign CPM[10379] = 12'b000000000000;
assign CPM[10380] = 12'b000000000000;
assign CPM[10381] = 12'b000000000000;
assign CPM[10382] = 12'b000000000000;
assign CPM[10383] = 12'b000000000000;
assign CPM[10384] = 12'b000000000000;
assign CPM[10385] = 12'b000000000000;
assign CPM[10386] = 12'b000000000000;
assign CPM[10387] = 12'b000000000000;
assign CPM[10388] = 12'b000000000000;
assign CPM[10389] = 12'b000000000000;
assign CPM[10390] = 12'b000000000000;
assign CPM[10391] = 12'b000000000000;
assign CPM[10392] = 12'b000000000000;
assign CPM[10393] = 12'b000000000000;
assign CPM[10394] = 12'b000000000000;
assign CPM[10395] = 12'b111111111111;
assign CPM[10396] = 12'b111111111111;
assign CPM[10397] = 12'b111111111111;
assign CPM[10398] = 12'b111111111111;
assign CPM[10399] = 12'b111111111111;
assign CPM[10400] = 12'b111111111111;
assign CPM[10401] = 12'b111111111111;
assign CPM[10402] = 12'b111111111111;
assign CPM[10403] = 12'b111111111111;
assign CPM[10404] = 12'b111111111111;
assign CPM[10405] = 12'b111111111111;
assign CPM[10406] = 12'b111111111111;
assign CPM[10407] = 12'b000000000000;
assign CPM[10408] = 12'b000000000000;
assign CPM[10409] = 12'b000000000000;
assign CPM[10410] = 12'b000000000000;
assign CPM[10411] = 12'b000000000000;
assign CPM[10412] = 12'b000000000000;
assign CPM[10413] = 12'b000000000000;
assign CPM[10414] = 12'b000000000000;
assign CPM[10415] = 12'b000000000000;
assign CPM[10416] = 12'b000000000000;
assign CPM[10417] = 12'b000000000000;
assign CPM[10418] = 12'b000000000000;
assign CPM[10419] = 12'b000000000000;
assign CPM[10420] = 12'b000000000000;
assign CPM[10421] = 12'b000000000000;
assign CPM[10422] = 12'b000000000000;
assign CPM[10423] = 12'b000000000000;
assign CPM[10424] = 12'b000000000000;
assign CPM[10425] = 12'b000000000000;
assign CPM[10426] = 12'b000000000000;
assign CPM[10427] = 12'b111111111111;
assign CPM[10428] = 12'b111111111111;
assign CPM[10429] = 12'b111111111111;
assign CPM[10430] = 12'b111111111111;
assign CPM[10431] = 12'b111111111111;
assign CPM[10432] = 12'b111111111111;
assign CPM[10433] = 12'b111111111111;
assign CPM[10434] = 12'b111111111111;
assign CPM[10435] = 12'b111111111111;
assign CPM[10436] = 12'b111111111111;
assign CPM[10437] = 12'b111111111111;
assign CPM[10438] = 12'b111111111111;
assign CPM[10439] = 12'b000000000000;
assign CPM[10440] = 12'b000000000000;
assign CPM[10441] = 12'b000000000000;
assign CPM[10442] = 12'b000000000000;
assign CPM[10443] = 12'b111111111111;
assign CPM[10444] = 12'b111111111111;
assign CPM[10445] = 12'b111111111111;
assign CPM[10446] = 12'b111111111111;
assign CPM[10447] = 12'b111111111111;
assign CPM[10448] = 12'b111111111111;
assign CPM[10449] = 12'b111111111111;
assign CPM[10450] = 12'b111111111111;
assign CPM[10451] = 12'b111111111111;
assign CPM[10452] = 12'b111111111111;
assign CPM[10453] = 12'b111111111111;
assign CPM[10454] = 12'b111111111111;
assign CPM[10455] = 12'b000000000000;
assign CPM[10456] = 12'b000000000000;
assign CPM[10457] = 12'b000000000000;
assign CPM[10458] = 12'b000000000000;
assign CPM[10459] = 12'b111111111111;
assign CPM[10460] = 12'b111111111111;
assign CPM[10461] = 12'b111111111111;
assign CPM[10462] = 12'b111111111111;
assign CPM[10463] = 12'b111111111111;
assign CPM[10464] = 12'b111111111111;
assign CPM[10465] = 12'b111111111111;
assign CPM[10466] = 12'b111111111111;
assign CPM[10467] = 12'b111111111111;
assign CPM[10468] = 12'b111111111111;
assign CPM[10469] = 12'b111111111111;
assign CPM[10470] = 12'b111111111111;
assign CPM[10471] = 12'b000000000000;
assign CPM[10472] = 12'b000000000000;
assign CPM[10473] = 12'b000000000000;
assign CPM[10474] = 12'b000000000000;
assign CPM[10475] = 12'b111111111111;
assign CPM[10476] = 12'b111111111111;
assign CPM[10477] = 12'b111111111111;
assign CPM[10478] = 12'b111111111111;
assign CPM[10479] = 12'b111111111111;
assign CPM[10480] = 12'b111111111111;
assign CPM[10481] = 12'b111111111111;
assign CPM[10482] = 12'b111111111111;
assign CPM[10483] = 12'b111111111111;
assign CPM[10484] = 12'b111111111111;
assign CPM[10485] = 12'b111111111111;
assign CPM[10486] = 12'b111111111111;
assign CPM[10487] = 12'b000000000000;
assign CPM[10488] = 12'b000000000000;
assign CPM[10489] = 12'b000000000000;
assign CPM[10490] = 12'b000000000000;
assign CPM[10491] = 12'b111111111111;
assign CPM[10492] = 12'b111111111111;
assign CPM[10493] = 12'b111111111111;
assign CPM[10494] = 12'b111111111111;
assign CPM[10495] = 12'b111111111111;
assign CPM[10496] = 12'b111111111111;
assign CPM[10497] = 12'b111111111111;
assign CPM[10498] = 12'b111111111111;
assign CPM[10499] = 12'b111111111111;
assign CPM[10500] = 12'b111111111111;
assign CPM[10501] = 12'b111111111111;
assign CPM[10502] = 12'b111111111111;
assign CPM[10503] = 12'b000000000000;
assign CPM[10504] = 12'b000000000000;
assign CPM[10505] = 12'b000000000000;
assign CPM[10506] = 12'b000000000000;
assign CPM[10507] = 12'b111111111111;
assign CPM[10508] = 12'b111111111111;
assign CPM[10509] = 12'b111111111111;
assign CPM[10510] = 12'b111111111111;
assign CPM[10511] = 12'b111111111111;
assign CPM[10512] = 12'b111111111111;
assign CPM[10513] = 12'b111111111111;
assign CPM[10514] = 12'b111111111111;
assign CPM[10515] = 12'b111111111111;
assign CPM[10516] = 12'b111111111111;
assign CPM[10517] = 12'b111111111111;
assign CPM[10518] = 12'b111111111111;
assign CPM[10519] = 12'b000000000000;
assign CPM[10520] = 12'b000000000000;
assign CPM[10521] = 12'b000000000000;
assign CPM[10522] = 12'b000000000000;
assign CPM[10523] = 12'b111111111111;
assign CPM[10524] = 12'b111111111111;
assign CPM[10525] = 12'b111111111111;
assign CPM[10526] = 12'b111111111111;
assign CPM[10527] = 12'b111111111111;
assign CPM[10528] = 12'b111111111111;
assign CPM[10529] = 12'b111111111111;
assign CPM[10530] = 12'b111111111111;
assign CPM[10531] = 12'b111111111111;
assign CPM[10532] = 12'b111111111111;
assign CPM[10533] = 12'b111111111111;
assign CPM[10534] = 12'b111111111111;
assign CPM[10535] = 12'b111111111111;
assign CPM[10536] = 12'b111111111111;
assign CPM[10537] = 12'b111111111111;
assign CPM[10538] = 12'b111111111111;
assign CPM[10539] = 12'b111111111111;
assign CPM[10540] = 12'b111111111111;
assign CPM[10541] = 12'b111111111111;
assign CPM[10542] = 12'b111111111111;
assign CPM[10543] = 12'b111111111111;
assign CPM[10544] = 12'b111111111111;
assign CPM[10545] = 12'b111111111111;
assign CPM[10546] = 12'b111111111111;
assign CPM[10547] = 12'b111111111111;
assign CPM[10548] = 12'b111111111111;
assign CPM[10549] = 12'b111111111111;
assign CPM[10550] = 12'b111111111111;
assign CPM[10551] = 12'b000000000000;
assign CPM[10552] = 12'b000000000000;
assign CPM[10553] = 12'b000000000000;
assign CPM[10554] = 12'b000000000000;
assign CPM[10555] = 12'b111111111111;
assign CPM[10556] = 12'b111111111111;
assign CPM[10557] = 12'b111111111111;
assign CPM[10558] = 12'b111111111111;
assign CPM[10559] = 12'b111111111111;
assign CPM[10560] = 12'b111111111111;
assign CPM[10561] = 12'b111111111111;
assign CPM[10562] = 12'b111111111111;
assign CPM[10563] = 12'b111111111111;
assign CPM[10564] = 12'b111111111111;
assign CPM[10565] = 12'b111111111111;
assign CPM[10566] = 12'b111111111111;
assign CPM[10567] = 12'b111111111111;
assign CPM[10568] = 12'b111111111111;
assign CPM[10569] = 12'b111111111111;
assign CPM[10570] = 12'b111111111111;
assign CPM[10571] = 12'b111111111111;
assign CPM[10572] = 12'b111111111111;
assign CPM[10573] = 12'b111111111111;
assign CPM[10574] = 12'b111111111111;
assign CPM[10575] = 12'b111111111111;
assign CPM[10576] = 12'b111111111111;
assign CPM[10577] = 12'b111111111111;
assign CPM[10578] = 12'b111111111111;
assign CPM[10579] = 12'b000000000000;
assign CPM[10580] = 12'b000000000000;
assign CPM[10581] = 12'b000000000000;
assign CPM[10582] = 12'b000000000000;
assign CPM[10583] = 12'b111111111111;
assign CPM[10584] = 12'b111111111111;
assign CPM[10585] = 12'b111111111111;
assign CPM[10586] = 12'b111111111111;
assign CPM[10587] = 12'b111111111111;
assign CPM[10588] = 12'b111111111111;
assign CPM[10589] = 12'b111111111111;
assign CPM[10590] = 12'b111111111111;
assign CPM[10591] = 12'b111111111111;
assign CPM[10592] = 12'b111111111111;
assign CPM[10593] = 12'b111111111111;
assign CPM[10594] = 12'b111111111111;
assign CPM[10595] = 12'b111111111111;
assign CPM[10596] = 12'b111111111111;
assign CPM[10597] = 12'b111111111111;
assign CPM[10598] = 12'b111111111111;
assign CPM[10599] = 12'b111111111111;
assign CPM[10600] = 12'b111111111111;
assign CPM[10601] = 12'b111111111111;
assign CPM[10602] = 12'b111111111111;
assign CPM[10603] = 12'b111111111111;
assign CPM[10604] = 12'b111111111111;
assign CPM[10605] = 12'b111111111111;
assign CPM[10606] = 12'b111111111111;
assign CPM[10607] = 12'b111111111111;
assign CPM[10608] = 12'b111111111111;
assign CPM[10609] = 12'b111111111111;
assign CPM[10610] = 12'b111111111111;
assign CPM[10611] = 12'b000000000000;
assign CPM[10612] = 12'b000000000000;
assign CPM[10613] = 12'b000000000000;
assign CPM[10614] = 12'b000000000000;
assign CPM[10615] = 12'b111111111111;
assign CPM[10616] = 12'b111111111111;
assign CPM[10617] = 12'b111111111111;
assign CPM[10618] = 12'b111111111111;
assign CPM[10619] = 12'b111111111111;
assign CPM[10620] = 12'b111111111111;
assign CPM[10621] = 12'b111111111111;
assign CPM[10622] = 12'b111111111111;
assign CPM[10623] = 12'b111111111111;
assign CPM[10624] = 12'b111111111111;
assign CPM[10625] = 12'b111111111111;
assign CPM[10626] = 12'b111111111111;
assign CPM[10627] = 12'b111111111111;
assign CPM[10628] = 12'b111111111111;
assign CPM[10629] = 12'b111111111111;
assign CPM[10630] = 12'b111111111111;
assign CPM[10631] = 12'b111111111111;
assign CPM[10632] = 12'b111111111111;
assign CPM[10633] = 12'b111111111111;
assign CPM[10634] = 12'b111111111111;
assign CPM[10635] = 12'b111111111111;
assign CPM[10636] = 12'b111111111111;
assign CPM[10637] = 12'b111111111111;
assign CPM[10638] = 12'b111111111111;
assign CPM[10639] = 12'b111111111111;
assign CPM[10640] = 12'b111111111111;
assign CPM[10641] = 12'b111111111111;
assign CPM[10642] = 12'b111111111111;
assign CPM[10643] = 12'b000000000000;
assign CPM[10644] = 12'b000000000000;
assign CPM[10645] = 12'b000000000000;
assign CPM[10646] = 12'b000000000000;
assign CPM[10647] = 12'b111111111111;
assign CPM[10648] = 12'b111111111111;
assign CPM[10649] = 12'b111111111111;
assign CPM[10650] = 12'b111111111111;
assign CPM[10651] = 12'b111111111111;
assign CPM[10652] = 12'b111111111111;
assign CPM[10653] = 12'b111111111111;
assign CPM[10654] = 12'b111111111111;
assign CPM[10655] = 12'b111111111111;
assign CPM[10656] = 12'b111111111111;
assign CPM[10657] = 12'b111111111111;
assign CPM[10658] = 12'b111111111111;
assign CPM[10659] = 12'b111111111111;
assign CPM[10660] = 12'b111111111111;
assign CPM[10661] = 12'b111111111111;
assign CPM[10662] = 12'b111111111111;
assign CPM[10663] = 12'b111111111111;
assign CPM[10664] = 12'b111111111111;
assign CPM[10665] = 12'b111111111111;
assign CPM[10666] = 12'b111111111111;
assign CPM[10667] = 12'b111111111111;
assign CPM[10668] = 12'b111111111111;
assign CPM[10669] = 12'b111111111111;
assign CPM[10670] = 12'b111111111111;
assign CPM[10671] = 12'b111111111111;
assign CPM[10672] = 12'b111111111111;
assign CPM[10673] = 12'b111111111111;
assign CPM[10674] = 12'b111111111111;
assign CPM[10675] = 12'b000000000000;
assign CPM[10676] = 12'b000000000000;
assign CPM[10677] = 12'b000000000000;
assign CPM[10678] = 12'b000000000000;
assign CPM[10679] = 12'b111111111111;
assign CPM[10680] = 12'b111111111111;
assign CPM[10681] = 12'b111111111111;
assign CPM[10682] = 12'b111111111111;
assign CPM[10683] = 12'b111111111111;
assign CPM[10684] = 12'b111111111111;
assign CPM[10685] = 12'b111111111111;
assign CPM[10686] = 12'b111111111111;
assign CPM[10687] = 12'b111111111111;
assign CPM[10688] = 12'b111111111111;
assign CPM[10689] = 12'b111111111111;
assign CPM[10690] = 12'b111111111111;
assign CPM[10691] = 12'b111111111111;
assign CPM[10692] = 12'b111111111111;
assign CPM[10693] = 12'b111111111111;
assign CPM[10694] = 12'b111111111111;
assign CPM[10695] = 12'b111111111111;
assign CPM[10696] = 12'b111111111111;
assign CPM[10697] = 12'b111111111111;
assign CPM[10698] = 12'b111111111111;
assign CPM[10699] = 12'b111111111111;
assign CPM[10700] = 12'b111111111111;
assign CPM[10701] = 12'b111111111111;
assign CPM[10702] = 12'b111111111111;
assign CPM[10703] = 12'b000000000000;
assign CPM[10704] = 12'b000000000000;
assign CPM[10705] = 12'b000000000000;
assign CPM[10706] = 12'b000000000000;
assign CPM[10707] = 12'b111111111111;
assign CPM[10708] = 12'b111111111111;
assign CPM[10709] = 12'b111111111111;
assign CPM[10710] = 12'b111111111111;
assign CPM[10711] = 12'b111111111111;
assign CPM[10712] = 12'b111111111111;
assign CPM[10713] = 12'b111111111111;
assign CPM[10714] = 12'b111111111111;
assign CPM[10715] = 12'b111111111111;
assign CPM[10716] = 12'b111111111111;
assign CPM[10717] = 12'b111111111111;
assign CPM[10718] = 12'b111111111111;
assign CPM[10719] = 12'b111111111111;
assign CPM[10720] = 12'b111111111111;
assign CPM[10721] = 12'b111111111111;
assign CPM[10722] = 12'b111111111111;
assign CPM[10723] = 12'b111111111111;
assign CPM[10724] = 12'b111111111111;
assign CPM[10725] = 12'b111111111111;
assign CPM[10726] = 12'b111111111111;
assign CPM[10727] = 12'b111111111111;
assign CPM[10728] = 12'b111111111111;
assign CPM[10729] = 12'b111111111111;
assign CPM[10730] = 12'b111111111111;
assign CPM[10731] = 12'b111111111111;
assign CPM[10732] = 12'b111111111111;
assign CPM[10733] = 12'b111111111111;
assign CPM[10734] = 12'b111111111111;
assign CPM[10735] = 12'b000000000000;
assign CPM[10736] = 12'b000000000000;
assign CPM[10737] = 12'b000000000000;
assign CPM[10738] = 12'b000000000000;
assign CPM[10739] = 12'b111111111111;
assign CPM[10740] = 12'b111111111111;
assign CPM[10741] = 12'b111111111111;
assign CPM[10742] = 12'b111111111111;
assign CPM[10743] = 12'b111111111111;
assign CPM[10744] = 12'b111111111111;
assign CPM[10745] = 12'b111111111111;
assign CPM[10746] = 12'b111111111111;
assign CPM[10747] = 12'b111111111111;
assign CPM[10748] = 12'b111111111111;
assign CPM[10749] = 12'b111111111111;
assign CPM[10750] = 12'b111111111111;
assign CPM[10751] = 12'b111111111111;
assign CPM[10752] = 12'b111111111111;
assign CPM[10753] = 12'b111111111111;
assign CPM[10754] = 12'b111111111111;
assign CPM[10755] = 12'b111111111111;
assign CPM[10756] = 12'b111111111111;
assign CPM[10757] = 12'b111111111111;
assign CPM[10758] = 12'b111111111111;
assign CPM[10759] = 12'b111111111111;
assign CPM[10760] = 12'b111111111111;
assign CPM[10761] = 12'b111111111111;
assign CPM[10762] = 12'b111111111111;
assign CPM[10763] = 12'b111111111111;
assign CPM[10764] = 12'b111111111111;
assign CPM[10765] = 12'b111111111111;
assign CPM[10766] = 12'b111111111111;
assign CPM[10767] = 12'b000000000000;
assign CPM[10768] = 12'b000000000000;
assign CPM[10769] = 12'b000000000000;
assign CPM[10770] = 12'b000000000000;
assign CPM[10771] = 12'b111111111111;
assign CPM[10772] = 12'b111111111111;
assign CPM[10773] = 12'b111111111111;
assign CPM[10774] = 12'b111111111111;
assign CPM[10775] = 12'b111111111111;
assign CPM[10776] = 12'b111111111111;
assign CPM[10777] = 12'b111111111111;
assign CPM[10778] = 12'b111111111111;
assign CPM[10779] = 12'b111111111111;
assign CPM[10780] = 12'b111111111111;
assign CPM[10781] = 12'b111111111111;
assign CPM[10782] = 12'b111111111111;
assign CPM[10783] = 12'b111111111111;
assign CPM[10784] = 12'b111111111111;
assign CPM[10785] = 12'b111111111111;
assign CPM[10786] = 12'b111111111111;
assign CPM[10787] = 12'b111111111111;
assign CPM[10788] = 12'b111111111111;
assign CPM[10789] = 12'b111111111111;
assign CPM[10790] = 12'b111111111111;
assign CPM[10791] = 12'b111111111111;
assign CPM[10792] = 12'b111111111111;
assign CPM[10793] = 12'b111111111111;
assign CPM[10794] = 12'b111111111111;
assign CPM[10795] = 12'b111111111111;
assign CPM[10796] = 12'b111111111111;
assign CPM[10797] = 12'b111111111111;
assign CPM[10798] = 12'b111111111111;
assign CPM[10799] = 12'b000000000000;
assign CPM[10800] = 12'b000000000000;
assign CPM[10801] = 12'b000000000000;
assign CPM[10802] = 12'b000000000000;
assign CPM[10803] = 12'b111111111111;
assign CPM[10804] = 12'b111111111111;
assign CPM[10805] = 12'b111111111111;
assign CPM[10806] = 12'b111111111111;
assign CPM[10807] = 12'b111111111111;
assign CPM[10808] = 12'b111111111111;
assign CPM[10809] = 12'b111111111111;
assign CPM[10810] = 12'b111111111111;
assign CPM[10811] = 12'b111111111111;
assign CPM[10812] = 12'b111111111111;
assign CPM[10813] = 12'b111111111111;
assign CPM[10814] = 12'b111111111111;
assign CPM[10815] = 12'b111111111111;
assign CPM[10816] = 12'b111111111111;
assign CPM[10817] = 12'b111111111111;
assign CPM[10818] = 12'b111111111111;
assign CPM[10819] = 12'b111111111111;
assign CPM[10820] = 12'b111111111111;
assign CPM[10821] = 12'b111111111111;
assign CPM[10822] = 12'b111111111111;
assign CPM[10823] = 12'b111111111111;
assign CPM[10824] = 12'b111111111111;
assign CPM[10825] = 12'b111111111111;
assign CPM[10826] = 12'b111111111111;
assign CPM[10827] = 12'b111111111111;
assign CPM[10828] = 12'b111111111111;
assign CPM[10829] = 12'b111111111111;
assign CPM[10830] = 12'b111111111111;
assign CPM[10831] = 12'b000000000000;
assign CPM[10832] = 12'b000000000000;
assign CPM[10833] = 12'b000000000000;
assign CPM[10834] = 12'b000000000000;
assign CPM[10835] = 12'b111111111111;
assign CPM[10836] = 12'b111111111111;
assign CPM[10837] = 12'b111111111111;
assign CPM[10838] = 12'b111111111111;
assign CPM[10839] = 12'b111111111111;
assign CPM[10840] = 12'b111111111111;
assign CPM[10841] = 12'b111111111111;
assign CPM[10842] = 12'b111111111111;
assign CPM[10843] = 12'b111111111111;
assign CPM[10844] = 12'b111111111111;
assign CPM[10845] = 12'b111111111111;
assign CPM[10846] = 12'b111111111111;
assign CPM[10847] = 12'b111111111111;
assign CPM[10848] = 12'b111111111111;
assign CPM[10849] = 12'b111111111111;
assign CPM[10850] = 12'b111111111111;
assign CPM[10851] = 12'b111111111111;
assign CPM[10852] = 12'b111111111111;
assign CPM[10853] = 12'b111111111111;
assign CPM[10854] = 12'b111111111111;
assign CPM[10855] = 12'b111111111111;
assign CPM[10856] = 12'b111111111111;
assign CPM[10857] = 12'b111111111111;
assign CPM[10858] = 12'b111111111111;
assign CPM[10859] = 12'b111111111111;
assign CPM[10860] = 12'b111111111111;
assign CPM[10861] = 12'b111111111111;
assign CPM[10862] = 12'b111111111111;
assign CPM[10863] = 12'b000000000000;
assign CPM[10864] = 12'b000000000000;
assign CPM[10865] = 12'b000000000000;
assign CPM[10866] = 12'b000000000000;
assign CPM[10867] = 12'b111111111111;
assign CPM[10868] = 12'b111111111111;
assign CPM[10869] = 12'b111111111111;
assign CPM[10870] = 12'b111111111111;
assign CPM[10871] = 12'b111111111111;
assign CPM[10872] = 12'b111111111111;
assign CPM[10873] = 12'b111111111111;
assign CPM[10874] = 12'b111111111111;
assign CPM[10875] = 12'b111111111111;
assign CPM[10876] = 12'b111111111111;
assign CPM[10877] = 12'b111111111111;
assign CPM[10878] = 12'b111111111111;
assign CPM[10879] = 12'b111111111111;
assign CPM[10880] = 12'b111111111111;
assign CPM[10881] = 12'b111111111111;
assign CPM[10882] = 12'b111111111111;
assign CPM[10883] = 12'b111111111111;
assign CPM[10884] = 12'b111111111111;
assign CPM[10885] = 12'b111111111111;
assign CPM[10886] = 12'b111111111111;
assign CPM[10887] = 12'b111111111111;
assign CPM[10888] = 12'b111111111111;
assign CPM[10889] = 12'b111111111111;
assign CPM[10890] = 12'b111111111111;
assign CPM[10891] = 12'b111111111111;
assign CPM[10892] = 12'b111111111111;
assign CPM[10893] = 12'b111111111111;
assign CPM[10894] = 12'b111111111111;
assign CPM[10895] = 12'b000000000000;
assign CPM[10896] = 12'b000000000000;
assign CPM[10897] = 12'b000000000000;
assign CPM[10898] = 12'b000000000000;
assign CPM[10899] = 12'b111111111111;
assign CPM[10900] = 12'b111111111111;
assign CPM[10901] = 12'b111111111111;
assign CPM[10902] = 12'b111111111111;
assign CPM[10903] = 12'b111111111111;
assign CPM[10904] = 12'b111111111111;
assign CPM[10905] = 12'b111111111111;
assign CPM[10906] = 12'b111111111111;
assign CPM[10907] = 12'b111111111111;
assign CPM[10908] = 12'b111111111111;
assign CPM[10909] = 12'b111111111111;
assign CPM[10910] = 12'b111111111111;
assign CPM[10911] = 12'b111111111111;
assign CPM[10912] = 12'b111111111111;
assign CPM[10913] = 12'b111111111111;
assign CPM[10914] = 12'b111111111111;
assign CPM[10915] = 12'b111111111111;
assign CPM[10916] = 12'b111111111111;
assign CPM[10917] = 12'b111111111111;
assign CPM[10918] = 12'b111111111111;
assign CPM[10919] = 12'b111111111111;
assign CPM[10920] = 12'b111111111111;
assign CPM[10921] = 12'b111111111111;
assign CPM[10922] = 12'b111111111111;
assign CPM[10923] = 12'b111111111111;
assign CPM[10924] = 12'b111111111111;
assign CPM[10925] = 12'b111111111111;
assign CPM[10926] = 12'b111111111111;
assign CPM[10927] = 12'b000000000000;
assign CPM[10928] = 12'b000000000000;
assign CPM[10929] = 12'b000000000000;
assign CPM[10930] = 12'b000000000000;
assign CPM[10931] = 12'b111111111111;
assign CPM[10932] = 12'b111111111111;
assign CPM[10933] = 12'b111111111111;
assign CPM[10934] = 12'b111111111111;
assign CPM[10935] = 12'b111111111111;
assign CPM[10936] = 12'b111111111111;
assign CPM[10937] = 12'b111111111111;
assign CPM[10938] = 12'b111111111111;
assign CPM[10939] = 12'b111111111111;
assign CPM[10940] = 12'b111111111111;
assign CPM[10941] = 12'b111111111111;
assign CPM[10942] = 12'b111111111111;
assign CPM[10943] = 12'b111111111111;
assign CPM[10944] = 12'b111111111111;
assign CPM[10945] = 12'b111111111111;
assign CPM[10946] = 12'b111111111111;
assign CPM[10947] = 12'b111111111111;
assign CPM[10948] = 12'b111111111111;
assign CPM[10949] = 12'b111111111111;
assign CPM[10950] = 12'b111111111111;
assign CPM[10951] = 12'b111111111111;
assign CPM[10952] = 12'b111111111111;
assign CPM[10953] = 12'b111111111111;
assign CPM[10954] = 12'b111111111111;
assign CPM[10955] = 12'b111111111111;
assign CPM[10956] = 12'b111111111111;
assign CPM[10957] = 12'b111111111111;
assign CPM[10958] = 12'b111111111111;
assign CPM[10959] = 12'b000000000000;
assign CPM[10960] = 12'b000000000000;
assign CPM[10961] = 12'b000000000000;
assign CPM[10962] = 12'b000000000000;
assign CPM[10963] = 12'b111111111111;
assign CPM[10964] = 12'b111111111111;
assign CPM[10965] = 12'b111111111111;
assign CPM[10966] = 12'b111111111111;
assign CPM[10967] = 12'b111111111111;
assign CPM[10968] = 12'b111111111111;
assign CPM[10969] = 12'b111111111111;
assign CPM[10970] = 12'b111111111111;
assign CPM[10971] = 12'b111111111111;
assign CPM[10972] = 12'b111111111111;
assign CPM[10973] = 12'b111111111111;
assign CPM[10974] = 12'b111111111111;
assign CPM[10975] = 12'b111111111111;
assign CPM[10976] = 12'b111111111111;
assign CPM[10977] = 12'b111111111111;
assign CPM[10978] = 12'b111111111111;
assign CPM[10979] = 12'b111111111111;
assign CPM[10980] = 12'b111111111111;
assign CPM[10981] = 12'b111111111111;
assign CPM[10982] = 12'b111111111111;
assign CPM[10983] = 12'b111111111111;
assign CPM[10984] = 12'b111111111111;
assign CPM[10985] = 12'b111111111111;
assign CPM[10986] = 12'b111111111111;
assign CPM[10987] = 12'b111111111111;
assign CPM[10988] = 12'b111111111111;
assign CPM[10989] = 12'b111111111111;
assign CPM[10990] = 12'b111111111111;
assign CPM[10991] = 12'b000000000000;
assign CPM[10992] = 12'b000000000000;
assign CPM[10993] = 12'b000000000000;
assign CPM[10994] = 12'b000000000000;
assign CPM[10995] = 12'b111111111111;
assign CPM[10996] = 12'b111111111111;
assign CPM[10997] = 12'b111111111111;
assign CPM[10998] = 12'b111111111111;
assign CPM[10999] = 12'b111111111111;
assign CPM[11000] = 12'b111111111111;
assign CPM[11001] = 12'b111111111111;
assign CPM[11002] = 12'b111111111111;
assign CPM[11003] = 12'b111111111111;
assign CPM[11004] = 12'b111111111111;
assign CPM[11005] = 12'b111111111111;
assign CPM[11006] = 12'b111111111111;
assign CPM[11007] = 12'b111111111111;
assign CPM[11008] = 12'b111111111111;
assign CPM[11009] = 12'b111111111111;
assign CPM[11010] = 12'b111111111111;
assign CPM[11011] = 12'b111111111111;
assign CPM[11012] = 12'b111111111111;
assign CPM[11013] = 12'b111111111111;
assign CPM[11014] = 12'b111111111111;
assign CPM[11015] = 12'b111111111111;
assign CPM[11016] = 12'b111111111111;
assign CPM[11017] = 12'b111111111111;
assign CPM[11018] = 12'b111111111111;
assign CPM[11019] = 12'b111111111111;
assign CPM[11020] = 12'b111111111111;
assign CPM[11021] = 12'b111111111111;
assign CPM[11022] = 12'b111111111111;
assign CPM[11023] = 12'b000000000000;
assign CPM[11024] = 12'b000000000000;
assign CPM[11025] = 12'b000000000000;
assign CPM[11026] = 12'b000000000000;
assign CPM[11027] = 12'b111111111111;
assign CPM[11028] = 12'b111111111111;
assign CPM[11029] = 12'b111111111111;
assign CPM[11030] = 12'b111111111111;
assign CPM[11031] = 12'b111111111111;
assign CPM[11032] = 12'b111111111111;
assign CPM[11033] = 12'b111111111111;
assign CPM[11034] = 12'b111111111111;
assign CPM[11035] = 12'b111111111111;
assign CPM[11036] = 12'b111111111111;
assign CPM[11037] = 12'b111111111111;
assign CPM[11038] = 12'b111111111111;
assign CPM[11039] = 12'b111111111111;
assign CPM[11040] = 12'b111111111111;
assign CPM[11041] = 12'b111111111111;
assign CPM[11042] = 12'b111111111111;
assign CPM[11043] = 12'b111111111111;
assign CPM[11044] = 12'b111111111111;
assign CPM[11045] = 12'b111111111111;
assign CPM[11046] = 12'b111111111111;
assign CPM[11047] = 12'b111111111111;
assign CPM[11048] = 12'b111111111111;
assign CPM[11049] = 12'b111111111111;
assign CPM[11050] = 12'b111111111111;
assign CPM[11051] = 12'b111111111111;
assign CPM[11052] = 12'b111111111111;
assign CPM[11053] = 12'b111111111111;
assign CPM[11054] = 12'b111111111111;
assign CPM[11055] = 12'b000000000000;
assign CPM[11056] = 12'b000000000000;
assign CPM[11057] = 12'b000000000000;
assign CPM[11058] = 12'b000000000000;
assign CPM[11059] = 12'b111111111111;
assign CPM[11060] = 12'b111111111111;
assign CPM[11061] = 12'b111111111111;
assign CPM[11062] = 12'b111111111111;
assign CPM[11063] = 12'b111111111111;
assign CPM[11064] = 12'b111111111111;
assign CPM[11065] = 12'b111111111111;
assign CPM[11066] = 12'b111111111111;
assign CPM[11067] = 12'b111111111111;
assign CPM[11068] = 12'b111111111111;
assign CPM[11069] = 12'b111111111111;
assign CPM[11070] = 12'b111111111111;
assign CPM[11071] = 12'b111111111111;
assign CPM[11072] = 12'b111111111111;
assign CPM[11073] = 12'b111111111111;
assign CPM[11074] = 12'b111111111111;
assign CPM[11075] = 12'b111111111111;
assign CPM[11076] = 12'b111111111111;
assign CPM[11077] = 12'b111111111111;
assign CPM[11078] = 12'b111111111111;
assign CPM[11079] = 12'b111111111111;
assign CPM[11080] = 12'b111111111111;
assign CPM[11081] = 12'b111111111111;
assign CPM[11082] = 12'b111111111111;
assign CPM[11083] = 12'b111111111111;
assign CPM[11084] = 12'b111111111111;
assign CPM[11085] = 12'b111111111111;
assign CPM[11086] = 12'b111111111111;
assign CPM[11087] = 12'b000000000000;
assign CPM[11088] = 12'b000000000000;
assign CPM[11089] = 12'b000000000000;
assign CPM[11090] = 12'b000000000000;
assign CPM[11091] = 12'b111111111111;
assign CPM[11092] = 12'b111111111111;
assign CPM[11093] = 12'b111111111111;
assign CPM[11094] = 12'b111111111111;
assign CPM[11095] = 12'b111111111111;
assign CPM[11096] = 12'b111111111111;
assign CPM[11097] = 12'b111111111111;
assign CPM[11098] = 12'b111111111111;
assign CPM[11099] = 12'b111111111111;
assign CPM[11100] = 12'b111111111111;
assign CPM[11101] = 12'b111111111111;
assign CPM[11102] = 12'b111111111111;
assign CPM[11103] = 12'b111111111111;
assign CPM[11104] = 12'b111111111111;
assign CPM[11105] = 12'b111111111111;
assign CPM[11106] = 12'b111111111111;
assign CPM[11107] = 12'b111111111111;
assign CPM[11108] = 12'b111111111111;
assign CPM[11109] = 12'b111111111111;
assign CPM[11110] = 12'b111111111111;
assign CPM[11111] = 12'b111111111111;
assign CPM[11112] = 12'b111111111111;
assign CPM[11113] = 12'b111111111111;
assign CPM[11114] = 12'b111111111111;
assign CPM[11115] = 12'b111111111111;
assign CPM[11116] = 12'b111111111111;
assign CPM[11117] = 12'b111111111111;
assign CPM[11118] = 12'b111111111111;
assign CPM[11119] = 12'b000000000000;
assign CPM[11120] = 12'b000000000000;
assign CPM[11121] = 12'b000000000000;
assign CPM[11122] = 12'b000000000000;
assign CPM[11123] = 12'b111111111111;
assign CPM[11124] = 12'b111111111111;
assign CPM[11125] = 12'b111111111111;
assign CPM[11126] = 12'b111111111111;
assign CPM[11127] = 12'b111111111111;
assign CPM[11128] = 12'b111111111111;
assign CPM[11129] = 12'b111111111111;
assign CPM[11130] = 12'b111111111111;
assign CPM[11131] = 12'b111111111111;
assign CPM[11132] = 12'b111111111111;
assign CPM[11133] = 12'b111111111111;
assign CPM[11134] = 12'b111111111111;
assign CPM[11135] = 12'b111111111111;
assign CPM[11136] = 12'b111111111111;
assign CPM[11137] = 12'b111111111111;
assign CPM[11138] = 12'b111111111111;
assign CPM[11139] = 12'b111111111111;
assign CPM[11140] = 12'b111111111111;
assign CPM[11141] = 12'b111111111111;
assign CPM[11142] = 12'b111111111111;
assign CPM[11143] = 12'b111111111111;
assign CPM[11144] = 12'b111111111111;
assign CPM[11145] = 12'b111111111111;
assign CPM[11146] = 12'b111111111111;
assign CPM[11147] = 12'b111111111111;
assign CPM[11148] = 12'b111111111111;
assign CPM[11149] = 12'b111111111111;
assign CPM[11150] = 12'b111111111111;
assign CPM[11151] = 12'b000000000000;
assign CPM[11152] = 12'b000000000000;
assign CPM[11153] = 12'b000000000000;
assign CPM[11154] = 12'b000000000000;
assign CPM[11155] = 12'b111111111111;
assign CPM[11156] = 12'b111111111111;
assign CPM[11157] = 12'b111111111111;
assign CPM[11158] = 12'b111111111111;
assign CPM[11159] = 12'b111111111111;
assign CPM[11160] = 12'b111111111111;
assign CPM[11161] = 12'b111111111111;
assign CPM[11162] = 12'b111111111111;
assign CPM[11163] = 12'b111111111111;
assign CPM[11164] = 12'b111111111111;
assign CPM[11165] = 12'b111111111111;
assign CPM[11166] = 12'b111111111111;
assign CPM[11167] = 12'b111111111111;
assign CPM[11168] = 12'b111111111111;
assign CPM[11169] = 12'b111111111111;
assign CPM[11170] = 12'b111111111111;
assign CPM[11171] = 12'b111111111111;
assign CPM[11172] = 12'b111111111111;
assign CPM[11173] = 12'b111111111111;
assign CPM[11174] = 12'b111111111111;
assign CPM[11175] = 12'b111111111111;
assign CPM[11176] = 12'b111111111111;
assign CPM[11177] = 12'b111111111111;
assign CPM[11178] = 12'b111111111111;
assign CPM[11179] = 12'b111111111111;
assign CPM[11180] = 12'b111111111111;
assign CPM[11181] = 12'b111111111111;
assign CPM[11182] = 12'b111111111111;
assign CPM[11183] = 12'b111111111111;
assign CPM[11184] = 12'b111111111111;
assign CPM[11185] = 12'b111111111111;
assign CPM[11186] = 12'b111111111111;
assign CPM[11187] = 12'b111111111111;
assign CPM[11188] = 12'b111111111111;
assign CPM[11189] = 12'b111111111111;
assign CPM[11190] = 12'b111111111111;
assign CPM[11191] = 12'b111111111111;
assign CPM[11192] = 12'b111111111111;
assign CPM[11193] = 12'b111111111111;
assign CPM[11194] = 12'b111111111111;
assign CPM[11195] = 12'b111111111111;
assign CPM[11196] = 12'b111111111111;
assign CPM[11197] = 12'b111111111111;
assign CPM[11198] = 12'b111111111111;
assign CPM[11199] = 12'b111111111111;
assign CPM[11200] = 12'b111111111111;
assign CPM[11201] = 12'b111111111111;
assign CPM[11202] = 12'b111111111111;
assign CPM[11203] = 12'b111111111111;
assign CPM[11204] = 12'b111111111111;
assign CPM[11205] = 12'b111111111111;
assign CPM[11206] = 12'b111111111111;
assign CPM[11207] = 12'b111111111111;
assign CPM[11208] = 12'b111111111111;
assign CPM[11209] = 12'b111111111111;
assign CPM[11210] = 12'b111111111111;
assign CPM[11211] = 12'b111111111111;
assign CPM[11212] = 12'b111111111111;
assign CPM[11213] = 12'b111111111111;
assign CPM[11214] = 12'b111111111111;
assign CPM[11215] = 12'b111111111111;
assign CPM[11216] = 12'b111111111111;
assign CPM[11217] = 12'b111111111111;
assign CPM[11218] = 12'b111111111111;
assign CPM[11219] = 12'b111111111111;
assign CPM[11220] = 12'b111111111111;
assign CPM[11221] = 12'b111111111111;
assign CPM[11222] = 12'b111111111111;
assign CPM[11223] = 12'b111111111111;
assign CPM[11224] = 12'b111111111111;
assign CPM[11225] = 12'b111111111111;
assign CPM[11226] = 12'b111111111111;
assign CPM[11227] = 12'b111111111111;
assign CPM[11228] = 12'b111111111111;
assign CPM[11229] = 12'b111111111111;
assign CPM[11230] = 12'b111111111111;
assign CPM[11231] = 12'b111111111111;
assign CPM[11232] = 12'b111111111111;
assign CPM[11233] = 12'b111111111111;
assign CPM[11234] = 12'b111111111111;
assign CPM[11235] = 12'b111111111111;
assign CPM[11236] = 12'b111111111111;
assign CPM[11237] = 12'b111111111111;
assign CPM[11238] = 12'b111111111111;
assign CPM[11239] = 12'b111111111111;
assign CPM[11240] = 12'b111111111111;
assign CPM[11241] = 12'b111111111111;
assign CPM[11242] = 12'b111111111111;
assign CPM[11243] = 12'b111111111111;
assign CPM[11244] = 12'b111111111111;
assign CPM[11245] = 12'b111111111111;
assign CPM[11246] = 12'b111111111111;
assign CPM[11247] = 12'b111111111111;
assign CPM[11248] = 12'b111111111111;
assign CPM[11249] = 12'b111111111111;
assign CPM[11250] = 12'b111111111111;
assign CPM[11251] = 12'b111111111111;
assign CPM[11252] = 12'b111111111111;
assign CPM[11253] = 12'b111111111111;
assign CPM[11254] = 12'b111111111111;
assign CPM[11255] = 12'b111111111111;
assign CPM[11256] = 12'b111111111111;
assign CPM[11257] = 12'b111111111111;
assign CPM[11258] = 12'b111111111111;
assign CPM[11259] = 12'b111111111111;
assign CPM[11260] = 12'b111111111111;
assign CPM[11261] = 12'b111111111111;
assign CPM[11262] = 12'b111111111111;
assign CPM[11263] = 12'b111111111111;
assign CPM[11264] = 12'b111111111111;
assign CPM[11265] = 12'b111111111111;
assign CPM[11266] = 12'b111111111111;
assign CPM[11267] = 12'b111111111111;
assign CPM[11268] = 12'b111111111111;
assign CPM[11269] = 12'b111111111111;
assign CPM[11270] = 12'b111111111111;
assign CPM[11271] = 12'b111111111111;
assign CPM[11272] = 12'b111111111111;
assign CPM[11273] = 12'b111111111111;
assign CPM[11274] = 12'b111111111111;
assign CPM[11275] = 12'b111111111111;
assign CPM[11276] = 12'b111111111111;
assign CPM[11277] = 12'b111111111111;
assign CPM[11278] = 12'b111111111111;
assign CPM[11279] = 12'b111111111111;
assign CPM[11280] = 12'b111111111111;
assign CPM[11281] = 12'b111111111111;
assign CPM[11282] = 12'b111111111111;
assign CPM[11283] = 12'b111111111111;
assign CPM[11284] = 12'b111111111111;
assign CPM[11285] = 12'b111111111111;
assign CPM[11286] = 12'b111111111111;
assign CPM[11287] = 12'b111111111111;
assign CPM[11288] = 12'b111111111111;
assign CPM[11289] = 12'b111111111111;
assign CPM[11290] = 12'b111111111111;
assign CPM[11291] = 12'b111111111111;
assign CPM[11292] = 12'b111111111111;
assign CPM[11293] = 12'b111111111111;
assign CPM[11294] = 12'b111111111111;
assign CPM[11295] = 12'b111111111111;
assign CPM[11296] = 12'b111111111111;
assign CPM[11297] = 12'b111111111111;
assign CPM[11298] = 12'b111111111111;
assign CPM[11299] = 12'b111111111111;
assign CPM[11300] = 12'b111111111111;
assign CPM[11301] = 12'b111111111111;
assign CPM[11302] = 12'b111111111111;
assign CPM[11303] = 12'b111111111111;
assign CPM[11304] = 12'b111111111111;
assign CPM[11305] = 12'b111111111111;
assign CPM[11306] = 12'b111111111111;
assign CPM[11307] = 12'b111111111111;
assign CPM[11308] = 12'b111111111111;
assign CPM[11309] = 12'b111111111111;
assign CPM[11310] = 12'b111111111111;
assign CPM[11311] = 12'b111111111111;
assign CPM[11312] = 12'b111111111111;
assign CPM[11313] = 12'b111111111111;
assign CPM[11314] = 12'b111111111111;
assign CPM[11315] = 12'b111111111111;
assign CPM[11316] = 12'b111111111111;
assign CPM[11317] = 12'b111111111111;
assign CPM[11318] = 12'b111111111111;
assign CPM[11319] = 12'b111111111111;
assign CPM[11320] = 12'b111111111111;
assign CPM[11321] = 12'b111111111111;
assign CPM[11322] = 12'b111111111111;
assign CPM[11323] = 12'b111111111111;
assign CPM[11324] = 12'b111111111111;
assign CPM[11325] = 12'b111111111111;
assign CPM[11326] = 12'b111111111111;
assign CPM[11327] = 12'b111111111111;
assign CPM[11328] = 12'b111111111111;
assign CPM[11329] = 12'b111111111111;
assign CPM[11330] = 12'b111111111111;
assign CPM[11331] = 12'b111111111111;
assign CPM[11332] = 12'b111111111111;
assign CPM[11333] = 12'b111111111111;
assign CPM[11334] = 12'b111111111111;
assign CPM[11335] = 12'b111111111111;
assign CPM[11336] = 12'b111111111111;
assign CPM[11337] = 12'b111111111111;
assign CPM[11338] = 12'b111111111111;
assign CPM[11339] = 12'b111111111111;
assign CPM[11340] = 12'b111111111111;
assign CPM[11341] = 12'b111111111111;
assign CPM[11342] = 12'b111111111111;
assign CPM[11343] = 12'b111111111111;
assign CPM[11344] = 12'b111111111111;
assign CPM[11345] = 12'b111111111111;
assign CPM[11346] = 12'b111111111111;
assign CPM[11347] = 12'b111111111111;
assign CPM[11348] = 12'b111111111111;
assign CPM[11349] = 12'b111111111111;
assign CPM[11350] = 12'b111111111111;
assign CPM[11351] = 12'b111111111111;
assign CPM[11352] = 12'b111111111111;
assign CPM[11353] = 12'b111111111111;
assign CPM[11354] = 12'b111111111111;
assign CPM[11355] = 12'b111111111111;
assign CPM[11356] = 12'b111111111111;
assign CPM[11357] = 12'b111111111111;
assign CPM[11358] = 12'b111111111111;
assign CPM[11359] = 12'b111111111111;
assign CPM[11360] = 12'b111111111111;
assign CPM[11361] = 12'b111111111111;
assign CPM[11362] = 12'b111111111111;
assign CPM[11363] = 12'b111111111111;
assign CPM[11364] = 12'b111111111111;
assign CPM[11365] = 12'b111111111111;
assign CPM[11366] = 12'b111111111111;
assign CPM[11367] = 12'b111111111111;
assign CPM[11368] = 12'b111111111111;
assign CPM[11369] = 12'b111111111111;
assign CPM[11370] = 12'b000000000000;
assign CPM[11371] = 12'b000000000000;
assign CPM[11372] = 12'b000000000000;
assign CPM[11373] = 12'b000000000000;
assign CPM[11374] = 12'b000000000000;
assign CPM[11375] = 12'b000000000000;
assign CPM[11376] = 12'b000000000000;
assign CPM[11377] = 12'b000000000000;
assign CPM[11378] = 12'b000000000000;
assign CPM[11379] = 12'b000000000000;
assign CPM[11380] = 12'b000000000000;
assign CPM[11381] = 12'b000000000000;
assign CPM[11382] = 12'b000000000000;
assign CPM[11383] = 12'b000000000000;
assign CPM[11384] = 12'b111111111111;
assign CPM[11385] = 12'b111111111111;
assign CPM[11386] = 12'b111111111111;
assign CPM[11387] = 12'b111111111111;
assign CPM[11388] = 12'b111111111111;
assign CPM[11389] = 12'b111111111111;
assign CPM[11390] = 12'b111111111111;
assign CPM[11391] = 12'b111111111111;
assign CPM[11392] = 12'b111111111111;
assign CPM[11393] = 12'b111111111111;
assign CPM[11394] = 12'b111111111111;
assign CPM[11395] = 12'b111111111111;
assign CPM[11396] = 12'b111111111111;
assign CPM[11397] = 12'b111111111111;
assign CPM[11398] = 12'b111111111111;
assign CPM[11399] = 12'b111111111111;
assign CPM[11400] = 12'b111111111111;
assign CPM[11401] = 12'b111111111111;
assign CPM[11402] = 12'b000000000000;
assign CPM[11403] = 12'b000000000000;
assign CPM[11404] = 12'b000000000000;
assign CPM[11405] = 12'b000000000000;
assign CPM[11406] = 12'b000000000000;
assign CPM[11407] = 12'b000000000000;
assign CPM[11408] = 12'b000000000000;
assign CPM[11409] = 12'b000000000000;
assign CPM[11410] = 12'b000000000000;
assign CPM[11411] = 12'b000000000000;
assign CPM[11412] = 12'b000000000000;
assign CPM[11413] = 12'b000000000000;
assign CPM[11414] = 12'b000000000000;
assign CPM[11415] = 12'b000000000000;
assign CPM[11416] = 12'b111111111111;
assign CPM[11417] = 12'b111111111111;
assign CPM[11418] = 12'b111111111111;
assign CPM[11419] = 12'b111111111111;
assign CPM[11420] = 12'b111111111111;
assign CPM[11421] = 12'b111111111111;
assign CPM[11422] = 12'b111111111111;
assign CPM[11423] = 12'b111111111111;
assign CPM[11424] = 12'b111111111111;
assign CPM[11425] = 12'b111111111111;
assign CPM[11426] = 12'b111111111111;
assign CPM[11427] = 12'b111111111111;
assign CPM[11428] = 12'b111111111111;
assign CPM[11429] = 12'b111111111111;
assign CPM[11430] = 12'b111111111111;
assign CPM[11431] = 12'b111111111111;
assign CPM[11432] = 12'b111111111111;
assign CPM[11433] = 12'b111111111111;
assign CPM[11434] = 12'b000000000000;
assign CPM[11435] = 12'b000000000000;
assign CPM[11436] = 12'b000000000000;
assign CPM[11437] = 12'b000000000000;
assign CPM[11438] = 12'b000000000000;
assign CPM[11439] = 12'b000000000000;
assign CPM[11440] = 12'b000000000000;
assign CPM[11441] = 12'b000000000000;
assign CPM[11442] = 12'b000000000000;
assign CPM[11443] = 12'b000000000000;
assign CPM[11444] = 12'b000000000000;
assign CPM[11445] = 12'b000000000000;
assign CPM[11446] = 12'b000000000000;
assign CPM[11447] = 12'b000000000000;
assign CPM[11448] = 12'b111111111111;
assign CPM[11449] = 12'b111111111111;
assign CPM[11450] = 12'b111111111111;
assign CPM[11451] = 12'b111111111111;
assign CPM[11452] = 12'b111111111111;
assign CPM[11453] = 12'b111111111111;
assign CPM[11454] = 12'b111111111111;
assign CPM[11455] = 12'b111111111111;
assign CPM[11456] = 12'b111111111111;
assign CPM[11457] = 12'b111111111111;
assign CPM[11458] = 12'b111111111111;
assign CPM[11459] = 12'b111111111111;
assign CPM[11460] = 12'b111111111111;
assign CPM[11461] = 12'b111111111111;
assign CPM[11462] = 12'b111111111111;
assign CPM[11463] = 12'b111111111111;
assign CPM[11464] = 12'b111111111111;
assign CPM[11465] = 12'b111111111111;
assign CPM[11466] = 12'b000000000000;
assign CPM[11467] = 12'b000000000000;
assign CPM[11468] = 12'b000000000000;
assign CPM[11469] = 12'b000000000000;
assign CPM[11470] = 12'b000000000000;
assign CPM[11471] = 12'b000000000000;
assign CPM[11472] = 12'b000000000000;
assign CPM[11473] = 12'b000000000000;
assign CPM[11474] = 12'b000000000000;
assign CPM[11475] = 12'b000000000000;
assign CPM[11476] = 12'b000000000000;
assign CPM[11477] = 12'b000000000000;
assign CPM[11478] = 12'b000000000000;
assign CPM[11479] = 12'b000000000000;
assign CPM[11480] = 12'b111111111111;
assign CPM[11481] = 12'b111111111111;
assign CPM[11482] = 12'b111111111111;
assign CPM[11483] = 12'b111111111111;
assign CPM[11484] = 12'b111111111111;
assign CPM[11485] = 12'b111111111111;
assign CPM[11486] = 12'b111111111111;
assign CPM[11487] = 12'b111111111111;
assign CPM[11488] = 12'b111111111111;
assign CPM[11489] = 12'b111111111111;
assign CPM[11490] = 12'b111111111111;
assign CPM[11491] = 12'b111111111111;
assign CPM[11492] = 12'b111111111111;
assign CPM[11493] = 12'b111111111111;
assign CPM[11494] = 12'b000000000000;
assign CPM[11495] = 12'b000000000000;
assign CPM[11496] = 12'b000000000000;
assign CPM[11497] = 12'b000000000000;
assign CPM[11498] = 12'b111111111111;
assign CPM[11499] = 12'b111111111111;
assign CPM[11500] = 12'b111111111111;
assign CPM[11501] = 12'b111111111111;
assign CPM[11502] = 12'b111111111111;
assign CPM[11503] = 12'b111111111111;
assign CPM[11504] = 12'b111111111111;
assign CPM[11505] = 12'b111111111111;
assign CPM[11506] = 12'b111111111111;
assign CPM[11507] = 12'b111111111111;
assign CPM[11508] = 12'b111111111111;
assign CPM[11509] = 12'b111111111111;
assign CPM[11510] = 12'b111111111111;
assign CPM[11511] = 12'b111111111111;
assign CPM[11512] = 12'b000000000000;
assign CPM[11513] = 12'b000000000000;
assign CPM[11514] = 12'b000000000000;
assign CPM[11515] = 12'b000000000000;
assign CPM[11516] = 12'b111111111111;
assign CPM[11517] = 12'b111111111111;
assign CPM[11518] = 12'b111111111111;
assign CPM[11519] = 12'b111111111111;
assign CPM[11520] = 12'b111111111111;
assign CPM[11521] = 12'b111111111111;
assign CPM[11522] = 12'b111111111111;
assign CPM[11523] = 12'b111111111111;
assign CPM[11524] = 12'b111111111111;
assign CPM[11525] = 12'b111111111111;
assign CPM[11526] = 12'b000000000000;
assign CPM[11527] = 12'b000000000000;
assign CPM[11528] = 12'b000000000000;
assign CPM[11529] = 12'b000000000000;
assign CPM[11530] = 12'b111111111111;
assign CPM[11531] = 12'b111111111111;
assign CPM[11532] = 12'b111111111111;
assign CPM[11533] = 12'b111111111111;
assign CPM[11534] = 12'b111111111111;
assign CPM[11535] = 12'b111111111111;
assign CPM[11536] = 12'b111111111111;
assign CPM[11537] = 12'b111111111111;
assign CPM[11538] = 12'b111111111111;
assign CPM[11539] = 12'b111111111111;
assign CPM[11540] = 12'b111111111111;
assign CPM[11541] = 12'b111111111111;
assign CPM[11542] = 12'b111111111111;
assign CPM[11543] = 12'b111111111111;
assign CPM[11544] = 12'b000000000000;
assign CPM[11545] = 12'b000000000000;
assign CPM[11546] = 12'b000000000000;
assign CPM[11547] = 12'b000000000000;
assign CPM[11548] = 12'b111111111111;
assign CPM[11549] = 12'b111111111111;
assign CPM[11550] = 12'b111111111111;
assign CPM[11551] = 12'b111111111111;
assign CPM[11552] = 12'b111111111111;
assign CPM[11553] = 12'b111111111111;
assign CPM[11554] = 12'b111111111111;
assign CPM[11555] = 12'b111111111111;
assign CPM[11556] = 12'b111111111111;
assign CPM[11557] = 12'b111111111111;
assign CPM[11558] = 12'b000000000000;
assign CPM[11559] = 12'b000000000000;
assign CPM[11560] = 12'b000000000000;
assign CPM[11561] = 12'b000000000000;
assign CPM[11562] = 12'b111111111111;
assign CPM[11563] = 12'b111111111111;
assign CPM[11564] = 12'b111111111111;
assign CPM[11565] = 12'b111111111111;
assign CPM[11566] = 12'b111111111111;
assign CPM[11567] = 12'b111111111111;
assign CPM[11568] = 12'b111111111111;
assign CPM[11569] = 12'b111111111111;
assign CPM[11570] = 12'b111111111111;
assign CPM[11571] = 12'b111111111111;
assign CPM[11572] = 12'b111111111111;
assign CPM[11573] = 12'b111111111111;
assign CPM[11574] = 12'b111111111111;
assign CPM[11575] = 12'b111111111111;
assign CPM[11576] = 12'b000000000000;
assign CPM[11577] = 12'b000000000000;
assign CPM[11578] = 12'b000000000000;
assign CPM[11579] = 12'b000000000000;
assign CPM[11580] = 12'b111111111111;
assign CPM[11581] = 12'b111111111111;
assign CPM[11582] = 12'b111111111111;
assign CPM[11583] = 12'b111111111111;
assign CPM[11584] = 12'b111111111111;
assign CPM[11585] = 12'b111111111111;
assign CPM[11586] = 12'b111111111111;
assign CPM[11587] = 12'b111111111111;
assign CPM[11588] = 12'b111111111111;
assign CPM[11589] = 12'b111111111111;
assign CPM[11590] = 12'b000000000000;
assign CPM[11591] = 12'b000000000000;
assign CPM[11592] = 12'b000000000000;
assign CPM[11593] = 12'b000000000000;
assign CPM[11594] = 12'b111111111111;
assign CPM[11595] = 12'b111111111111;
assign CPM[11596] = 12'b111111111111;
assign CPM[11597] = 12'b111111111111;
assign CPM[11598] = 12'b111111111111;
assign CPM[11599] = 12'b111111111111;
assign CPM[11600] = 12'b111111111111;
assign CPM[11601] = 12'b111111111111;
assign CPM[11602] = 12'b111111111111;
assign CPM[11603] = 12'b111111111111;
assign CPM[11604] = 12'b111111111111;
assign CPM[11605] = 12'b111111111111;
assign CPM[11606] = 12'b111111111111;
assign CPM[11607] = 12'b111111111111;
assign CPM[11608] = 12'b000000000000;
assign CPM[11609] = 12'b000000000000;
assign CPM[11610] = 12'b000000000000;
assign CPM[11611] = 12'b000000000000;
assign CPM[11612] = 12'b111111111111;
assign CPM[11613] = 12'b111111111111;
assign CPM[11614] = 12'b111111111111;
assign CPM[11615] = 12'b111111111111;
assign CPM[11616] = 12'b111111111111;
assign CPM[11617] = 12'b111111111111;
assign CPM[11618] = 12'b111111111111;
assign CPM[11619] = 12'b111111111111;
assign CPM[11620] = 12'b111111111111;
assign CPM[11621] = 12'b111111111111;
assign CPM[11622] = 12'b000000000000;
assign CPM[11623] = 12'b000000000000;
assign CPM[11624] = 12'b000000000000;
assign CPM[11625] = 12'b000000000000;
assign CPM[11626] = 12'b111111111111;
assign CPM[11627] = 12'b111111111111;
assign CPM[11628] = 12'b111111111111;
assign CPM[11629] = 12'b111111111111;
assign CPM[11630] = 12'b111111111111;
assign CPM[11631] = 12'b111111111111;
assign CPM[11632] = 12'b111111111111;
assign CPM[11633] = 12'b111111111111;
assign CPM[11634] = 12'b111111111111;
assign CPM[11635] = 12'b111111111111;
assign CPM[11636] = 12'b111111111111;
assign CPM[11637] = 12'b111111111111;
assign CPM[11638] = 12'b111111111111;
assign CPM[11639] = 12'b111111111111;
assign CPM[11640] = 12'b000000000000;
assign CPM[11641] = 12'b000000000000;
assign CPM[11642] = 12'b000000000000;
assign CPM[11643] = 12'b000000000000;
assign CPM[11644] = 12'b111111111111;
assign CPM[11645] = 12'b111111111111;
assign CPM[11646] = 12'b111111111111;
assign CPM[11647] = 12'b111111111111;
assign CPM[11648] = 12'b111111111111;
assign CPM[11649] = 12'b111111111111;
assign CPM[11650] = 12'b111111111111;
assign CPM[11651] = 12'b111111111111;
assign CPM[11652] = 12'b111111111111;
assign CPM[11653] = 12'b111111111111;
assign CPM[11654] = 12'b000000000000;
assign CPM[11655] = 12'b000000000000;
assign CPM[11656] = 12'b000000000000;
assign CPM[11657] = 12'b000000000000;
assign CPM[11658] = 12'b111111111111;
assign CPM[11659] = 12'b111111111111;
assign CPM[11660] = 12'b111111111111;
assign CPM[11661] = 12'b111111111111;
assign CPM[11662] = 12'b111111111111;
assign CPM[11663] = 12'b111111111111;
assign CPM[11664] = 12'b111111111111;
assign CPM[11665] = 12'b111111111111;
assign CPM[11666] = 12'b111111111111;
assign CPM[11667] = 12'b111111111111;
assign CPM[11668] = 12'b111111111111;
assign CPM[11669] = 12'b111111111111;
assign CPM[11670] = 12'b111111111111;
assign CPM[11671] = 12'b111111111111;
assign CPM[11672] = 12'b000000000000;
assign CPM[11673] = 12'b000000000000;
assign CPM[11674] = 12'b000000000000;
assign CPM[11675] = 12'b000000000000;
assign CPM[11676] = 12'b111111111111;
assign CPM[11677] = 12'b111111111111;
assign CPM[11678] = 12'b111111111111;
assign CPM[11679] = 12'b111111111111;
assign CPM[11680] = 12'b111111111111;
assign CPM[11681] = 12'b111111111111;
assign CPM[11682] = 12'b111111111111;
assign CPM[11683] = 12'b111111111111;
assign CPM[11684] = 12'b111111111111;
assign CPM[11685] = 12'b111111111111;
assign CPM[11686] = 12'b000000000000;
assign CPM[11687] = 12'b000000000000;
assign CPM[11688] = 12'b000000000000;
assign CPM[11689] = 12'b000000000000;
assign CPM[11690] = 12'b111111111111;
assign CPM[11691] = 12'b111111111111;
assign CPM[11692] = 12'b111111111111;
assign CPM[11693] = 12'b111111111111;
assign CPM[11694] = 12'b111111111111;
assign CPM[11695] = 12'b111111111111;
assign CPM[11696] = 12'b111111111111;
assign CPM[11697] = 12'b111111111111;
assign CPM[11698] = 12'b111111111111;
assign CPM[11699] = 12'b111111111111;
assign CPM[11700] = 12'b111111111111;
assign CPM[11701] = 12'b111111111111;
assign CPM[11702] = 12'b111111111111;
assign CPM[11703] = 12'b111111111111;
assign CPM[11704] = 12'b000000000000;
assign CPM[11705] = 12'b000000000000;
assign CPM[11706] = 12'b000000000000;
assign CPM[11707] = 12'b000000000000;
assign CPM[11708] = 12'b111111111111;
assign CPM[11709] = 12'b111111111111;
assign CPM[11710] = 12'b111111111111;
assign CPM[11711] = 12'b111111111111;
assign CPM[11712] = 12'b111111111111;
assign CPM[11713] = 12'b111111111111;
assign CPM[11714] = 12'b111111111111;
assign CPM[11715] = 12'b111111111111;
assign CPM[11716] = 12'b111111111111;
assign CPM[11717] = 12'b111111111111;
assign CPM[11718] = 12'b111111111111;
assign CPM[11719] = 12'b111111111111;
assign CPM[11720] = 12'b111111111111;
assign CPM[11721] = 12'b111111111111;
assign CPM[11722] = 12'b000000000000;
assign CPM[11723] = 12'b000000000000;
assign CPM[11724] = 12'b000000000000;
assign CPM[11725] = 12'b000000000000;
assign CPM[11726] = 12'b000000000000;
assign CPM[11727] = 12'b000000000000;
assign CPM[11728] = 12'b000000000000;
assign CPM[11729] = 12'b000000000000;
assign CPM[11730] = 12'b000000000000;
assign CPM[11731] = 12'b000000000000;
assign CPM[11732] = 12'b000000000000;
assign CPM[11733] = 12'b000000000000;
assign CPM[11734] = 12'b000000000000;
assign CPM[11735] = 12'b000000000000;
assign CPM[11736] = 12'b111111111111;
assign CPM[11737] = 12'b111111111111;
assign CPM[11738] = 12'b111111111111;
assign CPM[11739] = 12'b111111111111;
assign CPM[11740] = 12'b111111111111;
assign CPM[11741] = 12'b111111111111;
assign CPM[11742] = 12'b111111111111;
assign CPM[11743] = 12'b111111111111;
assign CPM[11744] = 12'b111111111111;
assign CPM[11745] = 12'b111111111111;
assign CPM[11746] = 12'b111111111111;
assign CPM[11747] = 12'b111111111111;
assign CPM[11748] = 12'b111111111111;
assign CPM[11749] = 12'b111111111111;
assign CPM[11750] = 12'b111111111111;
assign CPM[11751] = 12'b111111111111;
assign CPM[11752] = 12'b111111111111;
assign CPM[11753] = 12'b111111111111;
assign CPM[11754] = 12'b000000000000;
assign CPM[11755] = 12'b000000000000;
assign CPM[11756] = 12'b000000000000;
assign CPM[11757] = 12'b000000000000;
assign CPM[11758] = 12'b000000000000;
assign CPM[11759] = 12'b000000000000;
assign CPM[11760] = 12'b000000000000;
assign CPM[11761] = 12'b000000000000;
assign CPM[11762] = 12'b000000000000;
assign CPM[11763] = 12'b000000000000;
assign CPM[11764] = 12'b000000000000;
assign CPM[11765] = 12'b000000000000;
assign CPM[11766] = 12'b000000000000;
assign CPM[11767] = 12'b000000000000;
assign CPM[11768] = 12'b111111111111;
assign CPM[11769] = 12'b111111111111;
assign CPM[11770] = 12'b111111111111;
assign CPM[11771] = 12'b111111111111;
assign CPM[11772] = 12'b111111111111;
assign CPM[11773] = 12'b111111111111;
assign CPM[11774] = 12'b111111111111;
assign CPM[11775] = 12'b111111111111;
assign CPM[11776] = 12'b111111111111;
assign CPM[11777] = 12'b111111111111;
assign CPM[11778] = 12'b111111111111;
assign CPM[11779] = 12'b111111111111;
assign CPM[11780] = 12'b111111111111;
assign CPM[11781] = 12'b111111111111;
assign CPM[11782] = 12'b111111111111;
assign CPM[11783] = 12'b111111111111;
assign CPM[11784] = 12'b111111111111;
assign CPM[11785] = 12'b111111111111;
assign CPM[11786] = 12'b000000000000;
assign CPM[11787] = 12'b000000000000;
assign CPM[11788] = 12'b000000000000;
assign CPM[11789] = 12'b000000000000;
assign CPM[11790] = 12'b000000000000;
assign CPM[11791] = 12'b000000000000;
assign CPM[11792] = 12'b000000000000;
assign CPM[11793] = 12'b000000000000;
assign CPM[11794] = 12'b000000000000;
assign CPM[11795] = 12'b000000000000;
assign CPM[11796] = 12'b000000000000;
assign CPM[11797] = 12'b000000000000;
assign CPM[11798] = 12'b000000000000;
assign CPM[11799] = 12'b000000000000;
assign CPM[11800] = 12'b111111111111;
assign CPM[11801] = 12'b111111111111;
assign CPM[11802] = 12'b111111111111;
assign CPM[11803] = 12'b111111111111;
assign CPM[11804] = 12'b111111111111;
assign CPM[11805] = 12'b111111111111;
assign CPM[11806] = 12'b111111111111;
assign CPM[11807] = 12'b111111111111;
assign CPM[11808] = 12'b111111111111;
assign CPM[11809] = 12'b111111111111;
assign CPM[11810] = 12'b111111111111;
assign CPM[11811] = 12'b111111111111;
assign CPM[11812] = 12'b111111111111;
assign CPM[11813] = 12'b111111111111;
assign CPM[11814] = 12'b111111111111;
assign CPM[11815] = 12'b111111111111;
assign CPM[11816] = 12'b111111111111;
assign CPM[11817] = 12'b111111111111;
assign CPM[11818] = 12'b000000000000;
assign CPM[11819] = 12'b000000000000;
assign CPM[11820] = 12'b000000000000;
assign CPM[11821] = 12'b000000000000;
assign CPM[11822] = 12'b000000000000;
assign CPM[11823] = 12'b000000000000;
assign CPM[11824] = 12'b000000000000;
assign CPM[11825] = 12'b000000000000;
assign CPM[11826] = 12'b000000000000;
assign CPM[11827] = 12'b000000000000;
assign CPM[11828] = 12'b000000000000;
assign CPM[11829] = 12'b000000000000;
assign CPM[11830] = 12'b000000000000;
assign CPM[11831] = 12'b000000000000;
assign CPM[11832] = 12'b111111111111;
assign CPM[11833] = 12'b111111111111;
assign CPM[11834] = 12'b111111111111;
assign CPM[11835] = 12'b111111111111;
assign CPM[11836] = 12'b111111111111;
assign CPM[11837] = 12'b111111111111;
assign CPM[11838] = 12'b111111111111;
assign CPM[11839] = 12'b111111111111;
assign CPM[11840] = 12'b111111111111;
assign CPM[11841] = 12'b111111111111;
assign CPM[11842] = 12'b111111111111;
assign CPM[11843] = 12'b111111111111;
assign CPM[11844] = 12'b111111111111;
assign CPM[11845] = 12'b111111111111;
assign CPM[11846] = 12'b000000000000;
assign CPM[11847] = 12'b000000000000;
assign CPM[11848] = 12'b000000000000;
assign CPM[11849] = 12'b000000000000;
assign CPM[11850] = 12'b111111111111;
assign CPM[11851] = 12'b111111111111;
assign CPM[11852] = 12'b111111111111;
assign CPM[11853] = 12'b111111111111;
assign CPM[11854] = 12'b111111111111;
assign CPM[11855] = 12'b111111111111;
assign CPM[11856] = 12'b111111111111;
assign CPM[11857] = 12'b111111111111;
assign CPM[11858] = 12'b111111111111;
assign CPM[11859] = 12'b111111111111;
assign CPM[11860] = 12'b111111111111;
assign CPM[11861] = 12'b111111111111;
assign CPM[11862] = 12'b111111111111;
assign CPM[11863] = 12'b111111111111;
assign CPM[11864] = 12'b000000000000;
assign CPM[11865] = 12'b000000000000;
assign CPM[11866] = 12'b000000000000;
assign CPM[11867] = 12'b000000000000;
assign CPM[11868] = 12'b111111111111;
assign CPM[11869] = 12'b111111111111;
assign CPM[11870] = 12'b111111111111;
assign CPM[11871] = 12'b111111111111;
assign CPM[11872] = 12'b111111111111;
assign CPM[11873] = 12'b111111111111;
assign CPM[11874] = 12'b111111111111;
assign CPM[11875] = 12'b111111111111;
assign CPM[11876] = 12'b111111111111;
assign CPM[11877] = 12'b111111111111;
assign CPM[11878] = 12'b000000000000;
assign CPM[11879] = 12'b000000000000;
assign CPM[11880] = 12'b000000000000;
assign CPM[11881] = 12'b000000000000;
assign CPM[11882] = 12'b111111111111;
assign CPM[11883] = 12'b111111111111;
assign CPM[11884] = 12'b111111111111;
assign CPM[11885] = 12'b111111111111;
assign CPM[11886] = 12'b111111111111;
assign CPM[11887] = 12'b111111111111;
assign CPM[11888] = 12'b111111111111;
assign CPM[11889] = 12'b111111111111;
assign CPM[11890] = 12'b111111111111;
assign CPM[11891] = 12'b111111111111;
assign CPM[11892] = 12'b111111111111;
assign CPM[11893] = 12'b111111111111;
assign CPM[11894] = 12'b111111111111;
assign CPM[11895] = 12'b111111111111;
assign CPM[11896] = 12'b000000000000;
assign CPM[11897] = 12'b000000000000;
assign CPM[11898] = 12'b000000000000;
assign CPM[11899] = 12'b000000000000;
assign CPM[11900] = 12'b111111111111;
assign CPM[11901] = 12'b111111111111;
assign CPM[11902] = 12'b111111111111;
assign CPM[11903] = 12'b111111111111;
assign CPM[11904] = 12'b111111111111;
assign CPM[11905] = 12'b111111111111;
assign CPM[11906] = 12'b111111111111;
assign CPM[11907] = 12'b111111111111;
assign CPM[11908] = 12'b111111111111;
assign CPM[11909] = 12'b111111111111;
assign CPM[11910] = 12'b000000000000;
assign CPM[11911] = 12'b000000000000;
assign CPM[11912] = 12'b000000000000;
assign CPM[11913] = 12'b000000000000;
assign CPM[11914] = 12'b111111111111;
assign CPM[11915] = 12'b111111111111;
assign CPM[11916] = 12'b111111111111;
assign CPM[11917] = 12'b111111111111;
assign CPM[11918] = 12'b111111111111;
assign CPM[11919] = 12'b111111111111;
assign CPM[11920] = 12'b111111111111;
assign CPM[11921] = 12'b111111111111;
assign CPM[11922] = 12'b111111111111;
assign CPM[11923] = 12'b111111111111;
assign CPM[11924] = 12'b111111111111;
assign CPM[11925] = 12'b111111111111;
assign CPM[11926] = 12'b111111111111;
assign CPM[11927] = 12'b111111111111;
assign CPM[11928] = 12'b000000000000;
assign CPM[11929] = 12'b000000000000;
assign CPM[11930] = 12'b000000000000;
assign CPM[11931] = 12'b000000000000;
assign CPM[11932] = 12'b111111111111;
assign CPM[11933] = 12'b111111111111;
assign CPM[11934] = 12'b111111111111;
assign CPM[11935] = 12'b111111111111;
assign CPM[11936] = 12'b111111111111;
assign CPM[11937] = 12'b111111111111;
assign CPM[11938] = 12'b111111111111;
assign CPM[11939] = 12'b111111111111;
assign CPM[11940] = 12'b111111111111;
assign CPM[11941] = 12'b111111111111;
assign CPM[11942] = 12'b000000000000;
assign CPM[11943] = 12'b000000000000;
assign CPM[11944] = 12'b000000000000;
assign CPM[11945] = 12'b000000000000;
assign CPM[11946] = 12'b111111111111;
assign CPM[11947] = 12'b111111111111;
assign CPM[11948] = 12'b111111111111;
assign CPM[11949] = 12'b111111111111;
assign CPM[11950] = 12'b111111111111;
assign CPM[11951] = 12'b111111111111;
assign CPM[11952] = 12'b111111111111;
assign CPM[11953] = 12'b111111111111;
assign CPM[11954] = 12'b111111111111;
assign CPM[11955] = 12'b111111111111;
assign CPM[11956] = 12'b111111111111;
assign CPM[11957] = 12'b111111111111;
assign CPM[11958] = 12'b111111111111;
assign CPM[11959] = 12'b111111111111;
assign CPM[11960] = 12'b000000000000;
assign CPM[11961] = 12'b000000000000;
assign CPM[11962] = 12'b000000000000;
assign CPM[11963] = 12'b000000000000;
assign CPM[11964] = 12'b111111111111;
assign CPM[11965] = 12'b111111111111;
assign CPM[11966] = 12'b111111111111;
assign CPM[11967] = 12'b111111111111;
assign CPM[11968] = 12'b111111111111;
assign CPM[11969] = 12'b111111111111;
assign CPM[11970] = 12'b111111111111;
assign CPM[11971] = 12'b111111111111;
assign CPM[11972] = 12'b111111111111;
assign CPM[11973] = 12'b111111111111;
assign CPM[11974] = 12'b000000000000;
assign CPM[11975] = 12'b000000000000;
assign CPM[11976] = 12'b000000000000;
assign CPM[11977] = 12'b000000000000;
assign CPM[11978] = 12'b111111111111;
assign CPM[11979] = 12'b111111111111;
assign CPM[11980] = 12'b111111111111;
assign CPM[11981] = 12'b111111111111;
assign CPM[11982] = 12'b111111111111;
assign CPM[11983] = 12'b111111111111;
assign CPM[11984] = 12'b111111111111;
assign CPM[11985] = 12'b111111111111;
assign CPM[11986] = 12'b111111111111;
assign CPM[11987] = 12'b111111111111;
assign CPM[11988] = 12'b111111111111;
assign CPM[11989] = 12'b111111111111;
assign CPM[11990] = 12'b111111111111;
assign CPM[11991] = 12'b111111111111;
assign CPM[11992] = 12'b000000000000;
assign CPM[11993] = 12'b000000000000;
assign CPM[11994] = 12'b000000000000;
assign CPM[11995] = 12'b000000000000;
assign CPM[11996] = 12'b111111111111;
assign CPM[11997] = 12'b111111111111;
assign CPM[11998] = 12'b111111111111;
assign CPM[11999] = 12'b111111111111;
assign CPM[12000] = 12'b111111111111;
assign CPM[12001] = 12'b111111111111;
assign CPM[12002] = 12'b111111111111;
assign CPM[12003] = 12'b111111111111;
assign CPM[12004] = 12'b111111111111;
assign CPM[12005] = 12'b111111111111;
assign CPM[12006] = 12'b000000000000;
assign CPM[12007] = 12'b000000000000;
assign CPM[12008] = 12'b000000000000;
assign CPM[12009] = 12'b000000000000;
assign CPM[12010] = 12'b111111111111;
assign CPM[12011] = 12'b111111111111;
assign CPM[12012] = 12'b111111111111;
assign CPM[12013] = 12'b111111111111;
assign CPM[12014] = 12'b111111111111;
assign CPM[12015] = 12'b111111111111;
assign CPM[12016] = 12'b111111111111;
assign CPM[12017] = 12'b111111111111;
assign CPM[12018] = 12'b111111111111;
assign CPM[12019] = 12'b111111111111;
assign CPM[12020] = 12'b111111111111;
assign CPM[12021] = 12'b111111111111;
assign CPM[12022] = 12'b111111111111;
assign CPM[12023] = 12'b111111111111;
assign CPM[12024] = 12'b000000000000;
assign CPM[12025] = 12'b000000000000;
assign CPM[12026] = 12'b000000000000;
assign CPM[12027] = 12'b000000000000;
assign CPM[12028] = 12'b111111111111;
assign CPM[12029] = 12'b111111111111;
assign CPM[12030] = 12'b111111111111;
assign CPM[12031] = 12'b111111111111;
assign CPM[12032] = 12'b111111111111;
assign CPM[12033] = 12'b111111111111;
assign CPM[12034] = 12'b111111111111;
assign CPM[12035] = 12'b111111111111;
assign CPM[12036] = 12'b111111111111;
assign CPM[12037] = 12'b111111111111;
assign CPM[12038] = 12'b000000000000;
assign CPM[12039] = 12'b000000000000;
assign CPM[12040] = 12'b000000000000;
assign CPM[12041] = 12'b000000000000;
assign CPM[12042] = 12'b111111111111;
assign CPM[12043] = 12'b111111111111;
assign CPM[12044] = 12'b111111111111;
assign CPM[12045] = 12'b111111111111;
assign CPM[12046] = 12'b111111111111;
assign CPM[12047] = 12'b111111111111;
assign CPM[12048] = 12'b111111111111;
assign CPM[12049] = 12'b111111111111;
assign CPM[12050] = 12'b111111111111;
assign CPM[12051] = 12'b111111111111;
assign CPM[12052] = 12'b111111111111;
assign CPM[12053] = 12'b111111111111;
assign CPM[12054] = 12'b111111111111;
assign CPM[12055] = 12'b111111111111;
assign CPM[12056] = 12'b000000000000;
assign CPM[12057] = 12'b000000000000;
assign CPM[12058] = 12'b000000000000;
assign CPM[12059] = 12'b000000000000;
assign CPM[12060] = 12'b111111111111;
assign CPM[12061] = 12'b111111111111;
assign CPM[12062] = 12'b111111111111;
assign CPM[12063] = 12'b111111111111;
assign CPM[12064] = 12'b111111111111;
assign CPM[12065] = 12'b111111111111;
assign CPM[12066] = 12'b111111111111;
assign CPM[12067] = 12'b111111111111;
assign CPM[12068] = 12'b111111111111;
assign CPM[12069] = 12'b111111111111;
assign CPM[12070] = 12'b000000000000;
assign CPM[12071] = 12'b000000000000;
assign CPM[12072] = 12'b000000000000;
assign CPM[12073] = 12'b000000000000;
assign CPM[12074] = 12'b111111111111;
assign CPM[12075] = 12'b111111111111;
assign CPM[12076] = 12'b111111111111;
assign CPM[12077] = 12'b111111111111;
assign CPM[12078] = 12'b111111111111;
assign CPM[12079] = 12'b111111111111;
assign CPM[12080] = 12'b111111111111;
assign CPM[12081] = 12'b111111111111;
assign CPM[12082] = 12'b111111111111;
assign CPM[12083] = 12'b111111111111;
assign CPM[12084] = 12'b111111111111;
assign CPM[12085] = 12'b111111111111;
assign CPM[12086] = 12'b111111111111;
assign CPM[12087] = 12'b111111111111;
assign CPM[12088] = 12'b000000000000;
assign CPM[12089] = 12'b000000000000;
assign CPM[12090] = 12'b000000000000;
assign CPM[12091] = 12'b000000000000;
assign CPM[12092] = 12'b111111111111;
assign CPM[12093] = 12'b111111111111;
assign CPM[12094] = 12'b111111111111;
assign CPM[12095] = 12'b111111111111;
assign CPM[12096] = 12'b111111111111;
assign CPM[12097] = 12'b111111111111;
assign CPM[12098] = 12'b111111111111;
assign CPM[12099] = 12'b111111111111;
assign CPM[12100] = 12'b111111111111;
assign CPM[12101] = 12'b111111111111;
assign CPM[12102] = 12'b111111111111;
assign CPM[12103] = 12'b111111111111;
assign CPM[12104] = 12'b111111111111;
assign CPM[12105] = 12'b111111111111;
assign CPM[12106] = 12'b000000000000;
assign CPM[12107] = 12'b000000000000;
assign CPM[12108] = 12'b000000000000;
assign CPM[12109] = 12'b000000000000;
assign CPM[12110] = 12'b000000000000;
assign CPM[12111] = 12'b000000000000;
assign CPM[12112] = 12'b000000000000;
assign CPM[12113] = 12'b000000000000;
assign CPM[12114] = 12'b000000000000;
assign CPM[12115] = 12'b000000000000;
assign CPM[12116] = 12'b000000000000;
assign CPM[12117] = 12'b000000000000;
assign CPM[12118] = 12'b000000000000;
assign CPM[12119] = 12'b000000000000;
assign CPM[12120] = 12'b111111111111;
assign CPM[12121] = 12'b111111111111;
assign CPM[12122] = 12'b111111111111;
assign CPM[12123] = 12'b111111111111;
assign CPM[12124] = 12'b111111111111;
assign CPM[12125] = 12'b111111111111;
assign CPM[12126] = 12'b111111111111;
assign CPM[12127] = 12'b111111111111;
assign CPM[12128] = 12'b111111111111;
assign CPM[12129] = 12'b111111111111;
assign CPM[12130] = 12'b111111111111;
assign CPM[12131] = 12'b111111111111;
assign CPM[12132] = 12'b111111111111;
assign CPM[12133] = 12'b111111111111;
assign CPM[12134] = 12'b111111111111;
assign CPM[12135] = 12'b111111111111;
assign CPM[12136] = 12'b111111111111;
assign CPM[12137] = 12'b111111111111;
assign CPM[12138] = 12'b000000000000;
assign CPM[12139] = 12'b000000000000;
assign CPM[12140] = 12'b000000000000;
assign CPM[12141] = 12'b000000000000;
assign CPM[12142] = 12'b000000000000;
assign CPM[12143] = 12'b000000000000;
assign CPM[12144] = 12'b000000000000;
assign CPM[12145] = 12'b000000000000;
assign CPM[12146] = 12'b000000000000;
assign CPM[12147] = 12'b000000000000;
assign CPM[12148] = 12'b000000000000;
assign CPM[12149] = 12'b000000000000;
assign CPM[12150] = 12'b000000000000;
assign CPM[12151] = 12'b000000000000;
assign CPM[12152] = 12'b111111111111;
assign CPM[12153] = 12'b111111111111;
assign CPM[12154] = 12'b111111111111;
assign CPM[12155] = 12'b111111111111;
assign CPM[12156] = 12'b111111111111;
assign CPM[12157] = 12'b111111111111;
assign CPM[12158] = 12'b111111111111;
assign CPM[12159] = 12'b111111111111;
assign CPM[12160] = 12'b111111111111;
assign CPM[12161] = 12'b111111111111;
assign CPM[12162] = 12'b111111111111;
assign CPM[12163] = 12'b111111111111;
assign CPM[12164] = 12'b111111111111;
assign CPM[12165] = 12'b111111111111;
assign CPM[12166] = 12'b111111111111;
assign CPM[12167] = 12'b111111111111;
assign CPM[12168] = 12'b111111111111;
assign CPM[12169] = 12'b111111111111;
assign CPM[12170] = 12'b000000000000;
assign CPM[12171] = 12'b000000000000;
assign CPM[12172] = 12'b000000000000;
assign CPM[12173] = 12'b000000000000;
assign CPM[12174] = 12'b000000000000;
assign CPM[12175] = 12'b000000000000;
assign CPM[12176] = 12'b000000000000;
assign CPM[12177] = 12'b000000000000;
assign CPM[12178] = 12'b000000000000;
assign CPM[12179] = 12'b000000000000;
assign CPM[12180] = 12'b000000000000;
assign CPM[12181] = 12'b000000000000;
assign CPM[12182] = 12'b000000000000;
assign CPM[12183] = 12'b000000000000;
assign CPM[12184] = 12'b111111111111;
assign CPM[12185] = 12'b111111111111;
assign CPM[12186] = 12'b111111111111;
assign CPM[12187] = 12'b111111111111;
assign CPM[12188] = 12'b111111111111;
assign CPM[12189] = 12'b111111111111;
assign CPM[12190] = 12'b111111111111;
assign CPM[12191] = 12'b111111111111;
assign CPM[12192] = 12'b111111111111;
assign CPM[12193] = 12'b111111111111;
assign CPM[12194] = 12'b111111111111;
assign CPM[12195] = 12'b111111111111;
assign CPM[12196] = 12'b111111111111;
assign CPM[12197] = 12'b111111111111;
assign CPM[12198] = 12'b111111111111;
assign CPM[12199] = 12'b111111111111;
assign CPM[12200] = 12'b111111111111;
assign CPM[12201] = 12'b111111111111;
assign CPM[12202] = 12'b000000000000;
assign CPM[12203] = 12'b000000000000;
assign CPM[12204] = 12'b000000000000;
assign CPM[12205] = 12'b000000000000;
assign CPM[12206] = 12'b000000000000;
assign CPM[12207] = 12'b000000000000;
assign CPM[12208] = 12'b000000000000;
assign CPM[12209] = 12'b000000000000;
assign CPM[12210] = 12'b000000000000;
assign CPM[12211] = 12'b000000000000;
assign CPM[12212] = 12'b000000000000;
assign CPM[12213] = 12'b000000000000;
assign CPM[12214] = 12'b000000000000;
assign CPM[12215] = 12'b000000000000;
assign CPM[12216] = 12'b111111111111;
assign CPM[12217] = 12'b111111111111;
assign CPM[12218] = 12'b111111111111;
assign CPM[12219] = 12'b111111111111;
assign CPM[12220] = 12'b111111111111;
assign CPM[12221] = 12'b111111111111;
assign CPM[12222] = 12'b111111111111;
assign CPM[12223] = 12'b111111111111;
assign CPM[12224] = 12'b111111111111;
assign CPM[12225] = 12'b111111111111;
assign CPM[12226] = 12'b111111111111;
assign CPM[12227] = 12'b111111111111;
assign CPM[12228] = 12'b111111111111;
assign CPM[12229] = 12'b111111111111;
assign CPM[12230] = 12'b111111111111;
assign CPM[12231] = 12'b111111111111;
assign CPM[12232] = 12'b111111111111;
assign CPM[12233] = 12'b111111111111;
assign CPM[12234] = 12'b111111111111;
assign CPM[12235] = 12'b111111111111;
assign CPM[12236] = 12'b111111111111;
assign CPM[12237] = 12'b111111111111;
assign CPM[12238] = 12'b111111111111;
assign CPM[12239] = 12'b111111111111;
assign CPM[12240] = 12'b111111111111;
assign CPM[12241] = 12'b111111111111;
assign CPM[12242] = 12'b111111111111;
assign CPM[12243] = 12'b111111111111;
assign CPM[12244] = 12'b111111111111;
assign CPM[12245] = 12'b111111111111;
assign CPM[12246] = 12'b111111111111;
assign CPM[12247] = 12'b111111111111;
assign CPM[12248] = 12'b111111111111;
assign CPM[12249] = 12'b111111111111;
assign CPM[12250] = 12'b111111111111;
assign CPM[12251] = 12'b111111111111;
assign CPM[12252] = 12'b111111111111;
assign CPM[12253] = 12'b111111111111;
assign CPM[12254] = 12'b111111111111;
assign CPM[12255] = 12'b111111111111;
assign CPM[12256] = 12'b111111111111;
assign CPM[12257] = 12'b111111111111;
assign CPM[12258] = 12'b111111111111;
assign CPM[12259] = 12'b111111111111;
assign CPM[12260] = 12'b111111111111;
assign CPM[12261] = 12'b111111111111;
assign CPM[12262] = 12'b111111111111;
assign CPM[12263] = 12'b111111111111;
assign CPM[12264] = 12'b111111111111;
assign CPM[12265] = 12'b111111111111;
assign CPM[12266] = 12'b111111111111;
assign CPM[12267] = 12'b111111111111;
assign CPM[12268] = 12'b111111111111;
assign CPM[12269] = 12'b111111111111;
assign CPM[12270] = 12'b111111111111;
assign CPM[12271] = 12'b111111111111;
assign CPM[12272] = 12'b111111111111;
assign CPM[12273] = 12'b111111111111;
assign CPM[12274] = 12'b111111111111;
assign CPM[12275] = 12'b111111111111;
assign CPM[12276] = 12'b111111111111;
assign CPM[12277] = 12'b111111111111;
assign CPM[12278] = 12'b111111111111;
assign CPM[12279] = 12'b111111111111;
assign CPM[12280] = 12'b111111111111;
assign CPM[12281] = 12'b111111111111;
assign CPM[12282] = 12'b111111111111;
assign CPM[12283] = 12'b111111111111;
assign CPM[12284] = 12'b111111111111;
assign CPM[12285] = 12'b111111111111;
assign CPM[12286] = 12'b111111111111;
assign CPM[12287] = 12'b111111111111;
assign CPM[12288] = 12'b111111111111;
assign CPM[12289] = 12'b111111111111;
assign CPM[12290] = 12'b111111111111;
assign CPM[12291] = 12'b111111111111;
assign CPM[12292] = 12'b111111111111;
assign CPM[12293] = 12'b111111111111;
assign CPM[12294] = 12'b111111111111;
assign CPM[12295] = 12'b111111111111;
assign CPM[12296] = 12'b111111111111;
assign CPM[12297] = 12'b111111111111;
assign CPM[12298] = 12'b111111111111;
assign CPM[12299] = 12'b111111111111;
assign CPM[12300] = 12'b111111111111;
assign CPM[12301] = 12'b111111111111;
assign CPM[12302] = 12'b111111111111;
assign CPM[12303] = 12'b111111111111;
assign CPM[12304] = 12'b111111111111;
assign CPM[12305] = 12'b111111111111;
assign CPM[12306] = 12'b111111111111;
assign CPM[12307] = 12'b111111111111;
assign CPM[12308] = 12'b111111111111;
assign CPM[12309] = 12'b111111111111;
assign CPM[12310] = 12'b111111111111;
assign CPM[12311] = 12'b111111111111;
assign CPM[12312] = 12'b111111111111;
assign CPM[12313] = 12'b111111111111;
assign CPM[12314] = 12'b111111111111;
assign CPM[12315] = 12'b111111111111;
assign CPM[12316] = 12'b111111111111;
assign CPM[12317] = 12'b111111111111;
assign CPM[12318] = 12'b111111111111;
assign CPM[12319] = 12'b111111111111;
assign CPM[12320] = 12'b111111111111;
assign CPM[12321] = 12'b111111111111;
assign CPM[12322] = 12'b111111111111;
assign CPM[12323] = 12'b111111111111;
assign CPM[12324] = 12'b111111111111;
assign CPM[12325] = 12'b111111111111;
assign CPM[12326] = 12'b111111111111;
assign CPM[12327] = 12'b111111111111;
assign CPM[12328] = 12'b111111111111;
assign CPM[12329] = 12'b111111111111;
assign CPM[12330] = 12'b111111111111;
assign CPM[12331] = 12'b111111111111;
assign CPM[12332] = 12'b111111111111;
assign CPM[12333] = 12'b111111111111;
assign CPM[12334] = 12'b111111111111;
assign CPM[12335] = 12'b111111111111;
assign CPM[12336] = 12'b111111111111;
assign CPM[12337] = 12'b111111111111;
assign CPM[12338] = 12'b111111111111;
assign CPM[12339] = 12'b111111111111;
assign CPM[12340] = 12'b111111111111;
assign CPM[12341] = 12'b111111111111;
assign CPM[12342] = 12'b111111111111;
assign CPM[12343] = 12'b111111111111;
assign CPM[12344] = 12'b111111111111;
assign CPM[12345] = 12'b111111111111;
assign CPM[12346] = 12'b111111111111;
assign CPM[12347] = 12'b111111111111;
assign CPM[12348] = 12'b111111111111;
assign CPM[12349] = 12'b111111111111;
assign CPM[12350] = 12'b111111111111;
assign CPM[12351] = 12'b111111111111;
assign CPM[12352] = 12'b111111111111;
assign CPM[12353] = 12'b111111111111;
assign CPM[12354] = 12'b111111111111;
assign CPM[12355] = 12'b111111111111;
assign CPM[12356] = 12'b111111111111;
assign CPM[12357] = 12'b111111111111;
assign CPM[12358] = 12'b111111111111;
assign CPM[12359] = 12'b111111111111;
assign CPM[12360] = 12'b111111111111;
assign CPM[12361] = 12'b111111111111;
assign CPM[12362] = 12'b000000000000;
assign CPM[12363] = 12'b000000000000;
assign CPM[12364] = 12'b000000000000;
assign CPM[12365] = 12'b000000000000;
assign CPM[12366] = 12'b000000000000;
assign CPM[12367] = 12'b000000000000;
assign CPM[12368] = 12'b000000000000;
assign CPM[12369] = 12'b000000000000;
assign CPM[12370] = 12'b000000000000;
assign CPM[12371] = 12'b000000000000;
assign CPM[12372] = 12'b000000000000;
assign CPM[12373] = 12'b000000000000;
assign CPM[12374] = 12'b111111111111;
assign CPM[12375] = 12'b111111111111;
assign CPM[12376] = 12'b111111111111;
assign CPM[12377] = 12'b111111111111;
assign CPM[12378] = 12'b111111111111;
assign CPM[12379] = 12'b111111111111;
assign CPM[12380] = 12'b111111111111;
assign CPM[12381] = 12'b111111111111;
assign CPM[12382] = 12'b111111111111;
assign CPM[12383] = 12'b111111111111;
assign CPM[12384] = 12'b111111111111;
assign CPM[12385] = 12'b111111111111;
assign CPM[12386] = 12'b111111111111;
assign CPM[12387] = 12'b111111111111;
assign CPM[12388] = 12'b111111111111;
assign CPM[12389] = 12'b111111111111;
assign CPM[12390] = 12'b111111111111;
assign CPM[12391] = 12'b111111111111;
assign CPM[12392] = 12'b111111111111;
assign CPM[12393] = 12'b111111111111;
assign CPM[12394] = 12'b000000000000;
assign CPM[12395] = 12'b000000000000;
assign CPM[12396] = 12'b000000000000;
assign CPM[12397] = 12'b000000000000;
assign CPM[12398] = 12'b000000000000;
assign CPM[12399] = 12'b000000000000;
assign CPM[12400] = 12'b000000000000;
assign CPM[12401] = 12'b000000000000;
assign CPM[12402] = 12'b000000000000;
assign CPM[12403] = 12'b000000000000;
assign CPM[12404] = 12'b000000000000;
assign CPM[12405] = 12'b000000000000;
assign CPM[12406] = 12'b111111111111;
assign CPM[12407] = 12'b111111111111;
assign CPM[12408] = 12'b111111111111;
assign CPM[12409] = 12'b111111111111;
assign CPM[12410] = 12'b111111111111;
assign CPM[12411] = 12'b111111111111;
assign CPM[12412] = 12'b111111111111;
assign CPM[12413] = 12'b111111111111;
assign CPM[12414] = 12'b111111111111;
assign CPM[12415] = 12'b111111111111;
assign CPM[12416] = 12'b111111111111;
assign CPM[12417] = 12'b111111111111;
assign CPM[12418] = 12'b111111111111;
assign CPM[12419] = 12'b111111111111;
assign CPM[12420] = 12'b111111111111;
assign CPM[12421] = 12'b111111111111;
assign CPM[12422] = 12'b111111111111;
assign CPM[12423] = 12'b111111111111;
assign CPM[12424] = 12'b111111111111;
assign CPM[12425] = 12'b111111111111;
assign CPM[12426] = 12'b000000000000;
assign CPM[12427] = 12'b000000000000;
assign CPM[12428] = 12'b000000000000;
assign CPM[12429] = 12'b000000000000;
assign CPM[12430] = 12'b000000000000;
assign CPM[12431] = 12'b000000000000;
assign CPM[12432] = 12'b000000000000;
assign CPM[12433] = 12'b000000000000;
assign CPM[12434] = 12'b000000000000;
assign CPM[12435] = 12'b000000000000;
assign CPM[12436] = 12'b000000000000;
assign CPM[12437] = 12'b000000000000;
assign CPM[12438] = 12'b111111111111;
assign CPM[12439] = 12'b111111111111;
assign CPM[12440] = 12'b111111111111;
assign CPM[12441] = 12'b111111111111;
assign CPM[12442] = 12'b111111111111;
assign CPM[12443] = 12'b111111111111;
assign CPM[12444] = 12'b111111111111;
assign CPM[12445] = 12'b111111111111;
assign CPM[12446] = 12'b111111111111;
assign CPM[12447] = 12'b111111111111;
assign CPM[12448] = 12'b111111111111;
assign CPM[12449] = 12'b111111111111;
assign CPM[12450] = 12'b111111111111;
assign CPM[12451] = 12'b111111111111;
assign CPM[12452] = 12'b111111111111;
assign CPM[12453] = 12'b111111111111;
assign CPM[12454] = 12'b111111111111;
assign CPM[12455] = 12'b111111111111;
assign CPM[12456] = 12'b111111111111;
assign CPM[12457] = 12'b111111111111;
assign CPM[12458] = 12'b000000000000;
assign CPM[12459] = 12'b000000000000;
assign CPM[12460] = 12'b000000000000;
assign CPM[12461] = 12'b000000000000;
assign CPM[12462] = 12'b000000000000;
assign CPM[12463] = 12'b000000000000;
assign CPM[12464] = 12'b000000000000;
assign CPM[12465] = 12'b000000000000;
assign CPM[12466] = 12'b000000000000;
assign CPM[12467] = 12'b000000000000;
assign CPM[12468] = 12'b000000000000;
assign CPM[12469] = 12'b000000000000;
assign CPM[12470] = 12'b111111111111;
assign CPM[12471] = 12'b111111111111;
assign CPM[12472] = 12'b111111111111;
assign CPM[12473] = 12'b111111111111;
assign CPM[12474] = 12'b111111111111;
assign CPM[12475] = 12'b111111111111;
assign CPM[12476] = 12'b111111111111;
assign CPM[12477] = 12'b111111111111;
assign CPM[12478] = 12'b111111111111;
assign CPM[12479] = 12'b111111111111;
assign CPM[12480] = 12'b111111111111;
assign CPM[12481] = 12'b111111111111;
assign CPM[12482] = 12'b111111111111;
assign CPM[12483] = 12'b111111111111;
assign CPM[12484] = 12'b111111111111;
assign CPM[12485] = 12'b111111111111;
assign CPM[12486] = 12'b000000000000;
assign CPM[12487] = 12'b000000000000;
assign CPM[12488] = 12'b000000000000;
assign CPM[12489] = 12'b000000000000;
assign CPM[12490] = 12'b111111111111;
assign CPM[12491] = 12'b111111111111;
assign CPM[12492] = 12'b111111111111;
assign CPM[12493] = 12'b111111111111;
assign CPM[12494] = 12'b111111111111;
assign CPM[12495] = 12'b111111111111;
assign CPM[12496] = 12'b111111111111;
assign CPM[12497] = 12'b111111111111;
assign CPM[12498] = 12'b111111111111;
assign CPM[12499] = 12'b111111111111;
assign CPM[12500] = 12'b111111111111;
assign CPM[12501] = 12'b111111111111;
assign CPM[12502] = 12'b000000000000;
assign CPM[12503] = 12'b000000000000;
assign CPM[12504] = 12'b000000000000;
assign CPM[12505] = 12'b000000000000;
assign CPM[12506] = 12'b111111111111;
assign CPM[12507] = 12'b111111111111;
assign CPM[12508] = 12'b111111111111;
assign CPM[12509] = 12'b111111111111;
assign CPM[12510] = 12'b111111111111;
assign CPM[12511] = 12'b111111111111;
assign CPM[12512] = 12'b111111111111;
assign CPM[12513] = 12'b111111111111;
assign CPM[12514] = 12'b111111111111;
assign CPM[12515] = 12'b111111111111;
assign CPM[12516] = 12'b111111111111;
assign CPM[12517] = 12'b111111111111;
assign CPM[12518] = 12'b000000000000;
assign CPM[12519] = 12'b000000000000;
assign CPM[12520] = 12'b000000000000;
assign CPM[12521] = 12'b000000000000;
assign CPM[12522] = 12'b111111111111;
assign CPM[12523] = 12'b111111111111;
assign CPM[12524] = 12'b111111111111;
assign CPM[12525] = 12'b111111111111;
assign CPM[12526] = 12'b111111111111;
assign CPM[12527] = 12'b111111111111;
assign CPM[12528] = 12'b111111111111;
assign CPM[12529] = 12'b111111111111;
assign CPM[12530] = 12'b111111111111;
assign CPM[12531] = 12'b111111111111;
assign CPM[12532] = 12'b111111111111;
assign CPM[12533] = 12'b111111111111;
assign CPM[12534] = 12'b000000000000;
assign CPM[12535] = 12'b000000000000;
assign CPM[12536] = 12'b000000000000;
assign CPM[12537] = 12'b000000000000;
assign CPM[12538] = 12'b111111111111;
assign CPM[12539] = 12'b111111111111;
assign CPM[12540] = 12'b111111111111;
assign CPM[12541] = 12'b111111111111;
assign CPM[12542] = 12'b111111111111;
assign CPM[12543] = 12'b111111111111;
assign CPM[12544] = 12'b111111111111;
assign CPM[12545] = 12'b111111111111;
assign CPM[12546] = 12'b111111111111;
assign CPM[12547] = 12'b111111111111;
assign CPM[12548] = 12'b111111111111;
assign CPM[12549] = 12'b111111111111;
assign CPM[12550] = 12'b000000000000;
assign CPM[12551] = 12'b000000000000;
assign CPM[12552] = 12'b000000000000;
assign CPM[12553] = 12'b000000000000;
assign CPM[12554] = 12'b111111111111;
assign CPM[12555] = 12'b111111111111;
assign CPM[12556] = 12'b111111111111;
assign CPM[12557] = 12'b111111111111;
assign CPM[12558] = 12'b111111111111;
assign CPM[12559] = 12'b111111111111;
assign CPM[12560] = 12'b111111111111;
assign CPM[12561] = 12'b111111111111;
assign CPM[12562] = 12'b111111111111;
assign CPM[12563] = 12'b111111111111;
assign CPM[12564] = 12'b111111111111;
assign CPM[12565] = 12'b111111111111;
assign CPM[12566] = 12'b000000000000;
assign CPM[12567] = 12'b000000000000;
assign CPM[12568] = 12'b000000000000;
assign CPM[12569] = 12'b000000000000;
assign CPM[12570] = 12'b111111111111;
assign CPM[12571] = 12'b111111111111;
assign CPM[12572] = 12'b111111111111;
assign CPM[12573] = 12'b111111111111;
assign CPM[12574] = 12'b111111111111;
assign CPM[12575] = 12'b111111111111;
assign CPM[12576] = 12'b111111111111;
assign CPM[12577] = 12'b111111111111;
assign CPM[12578] = 12'b111111111111;
assign CPM[12579] = 12'b111111111111;
assign CPM[12580] = 12'b111111111111;
assign CPM[12581] = 12'b111111111111;
assign CPM[12582] = 12'b000000000000;
assign CPM[12583] = 12'b000000000000;
assign CPM[12584] = 12'b000000000000;
assign CPM[12585] = 12'b000000000000;
assign CPM[12586] = 12'b111111111111;
assign CPM[12587] = 12'b111111111111;
assign CPM[12588] = 12'b111111111111;
assign CPM[12589] = 12'b111111111111;
assign CPM[12590] = 12'b111111111111;
assign CPM[12591] = 12'b111111111111;
assign CPM[12592] = 12'b111111111111;
assign CPM[12593] = 12'b111111111111;
assign CPM[12594] = 12'b111111111111;
assign CPM[12595] = 12'b111111111111;
assign CPM[12596] = 12'b111111111111;
assign CPM[12597] = 12'b111111111111;
assign CPM[12598] = 12'b000000000000;
assign CPM[12599] = 12'b000000000000;
assign CPM[12600] = 12'b000000000000;
assign CPM[12601] = 12'b000000000000;
assign CPM[12602] = 12'b111111111111;
assign CPM[12603] = 12'b111111111111;
assign CPM[12604] = 12'b111111111111;
assign CPM[12605] = 12'b111111111111;
assign CPM[12606] = 12'b111111111111;
assign CPM[12607] = 12'b111111111111;
assign CPM[12608] = 12'b111111111111;
assign CPM[12609] = 12'b111111111111;
assign CPM[12610] = 12'b111111111111;
assign CPM[12611] = 12'b111111111111;
assign CPM[12612] = 12'b111111111111;
assign CPM[12613] = 12'b111111111111;
assign CPM[12614] = 12'b000000000000;
assign CPM[12615] = 12'b000000000000;
assign CPM[12616] = 12'b000000000000;
assign CPM[12617] = 12'b000000000000;
assign CPM[12618] = 12'b111111111111;
assign CPM[12619] = 12'b111111111111;
assign CPM[12620] = 12'b111111111111;
assign CPM[12621] = 12'b111111111111;
assign CPM[12622] = 12'b111111111111;
assign CPM[12623] = 12'b111111111111;
assign CPM[12624] = 12'b111111111111;
assign CPM[12625] = 12'b111111111111;
assign CPM[12626] = 12'b111111111111;
assign CPM[12627] = 12'b111111111111;
assign CPM[12628] = 12'b111111111111;
assign CPM[12629] = 12'b111111111111;
assign CPM[12630] = 12'b000000000000;
assign CPM[12631] = 12'b000000000000;
assign CPM[12632] = 12'b000000000000;
assign CPM[12633] = 12'b000000000000;
assign CPM[12634] = 12'b111111111111;
assign CPM[12635] = 12'b111111111111;
assign CPM[12636] = 12'b111111111111;
assign CPM[12637] = 12'b111111111111;
assign CPM[12638] = 12'b111111111111;
assign CPM[12639] = 12'b111111111111;
assign CPM[12640] = 12'b111111111111;
assign CPM[12641] = 12'b111111111111;
assign CPM[12642] = 12'b111111111111;
assign CPM[12643] = 12'b111111111111;
assign CPM[12644] = 12'b111111111111;
assign CPM[12645] = 12'b111111111111;
assign CPM[12646] = 12'b000000000000;
assign CPM[12647] = 12'b000000000000;
assign CPM[12648] = 12'b000000000000;
assign CPM[12649] = 12'b000000000000;
assign CPM[12650] = 12'b111111111111;
assign CPM[12651] = 12'b111111111111;
assign CPM[12652] = 12'b111111111111;
assign CPM[12653] = 12'b111111111111;
assign CPM[12654] = 12'b111111111111;
assign CPM[12655] = 12'b111111111111;
assign CPM[12656] = 12'b111111111111;
assign CPM[12657] = 12'b111111111111;
assign CPM[12658] = 12'b111111111111;
assign CPM[12659] = 12'b111111111111;
assign CPM[12660] = 12'b111111111111;
assign CPM[12661] = 12'b111111111111;
assign CPM[12662] = 12'b000000000000;
assign CPM[12663] = 12'b000000000000;
assign CPM[12664] = 12'b000000000000;
assign CPM[12665] = 12'b000000000000;
assign CPM[12666] = 12'b111111111111;
assign CPM[12667] = 12'b111111111111;
assign CPM[12668] = 12'b111111111111;
assign CPM[12669] = 12'b111111111111;
assign CPM[12670] = 12'b111111111111;
assign CPM[12671] = 12'b111111111111;
assign CPM[12672] = 12'b111111111111;
assign CPM[12673] = 12'b111111111111;
assign CPM[12674] = 12'b111111111111;
assign CPM[12675] = 12'b111111111111;
assign CPM[12676] = 12'b111111111111;
assign CPM[12677] = 12'b111111111111;
assign CPM[12678] = 12'b000000000000;
assign CPM[12679] = 12'b000000000000;
assign CPM[12680] = 12'b000000000000;
assign CPM[12681] = 12'b000000000000;
assign CPM[12682] = 12'b111111111111;
assign CPM[12683] = 12'b111111111111;
assign CPM[12684] = 12'b111111111111;
assign CPM[12685] = 12'b111111111111;
assign CPM[12686] = 12'b111111111111;
assign CPM[12687] = 12'b111111111111;
assign CPM[12688] = 12'b111111111111;
assign CPM[12689] = 12'b111111111111;
assign CPM[12690] = 12'b111111111111;
assign CPM[12691] = 12'b111111111111;
assign CPM[12692] = 12'b111111111111;
assign CPM[12693] = 12'b111111111111;
assign CPM[12694] = 12'b000000000000;
assign CPM[12695] = 12'b000000000000;
assign CPM[12696] = 12'b000000000000;
assign CPM[12697] = 12'b000000000000;
assign CPM[12698] = 12'b111111111111;
assign CPM[12699] = 12'b111111111111;
assign CPM[12700] = 12'b111111111111;
assign CPM[12701] = 12'b111111111111;
assign CPM[12702] = 12'b111111111111;
assign CPM[12703] = 12'b111111111111;
assign CPM[12704] = 12'b111111111111;
assign CPM[12705] = 12'b111111111111;
assign CPM[12706] = 12'b111111111111;
assign CPM[12707] = 12'b111111111111;
assign CPM[12708] = 12'b111111111111;
assign CPM[12709] = 12'b111111111111;
assign CPM[12710] = 12'b111111111111;
assign CPM[12711] = 12'b111111111111;
assign CPM[12712] = 12'b111111111111;
assign CPM[12713] = 12'b111111111111;
assign CPM[12714] = 12'b000000000000;
assign CPM[12715] = 12'b000000000000;
assign CPM[12716] = 12'b000000000000;
assign CPM[12717] = 12'b000000000000;
assign CPM[12718] = 12'b000000000000;
assign CPM[12719] = 12'b000000000000;
assign CPM[12720] = 12'b000000000000;
assign CPM[12721] = 12'b000000000000;
assign CPM[12722] = 12'b000000000000;
assign CPM[12723] = 12'b000000000000;
assign CPM[12724] = 12'b000000000000;
assign CPM[12725] = 12'b000000000000;
assign CPM[12726] = 12'b000000000000;
assign CPM[12727] = 12'b000000000000;
assign CPM[12728] = 12'b000000000000;
assign CPM[12729] = 12'b000000000000;
assign CPM[12730] = 12'b111111111111;
assign CPM[12731] = 12'b111111111111;
assign CPM[12732] = 12'b111111111111;
assign CPM[12733] = 12'b111111111111;
assign CPM[12734] = 12'b111111111111;
assign CPM[12735] = 12'b111111111111;
assign CPM[12736] = 12'b111111111111;
assign CPM[12737] = 12'b111111111111;
assign CPM[12738] = 12'b111111111111;
assign CPM[12739] = 12'b111111111111;
assign CPM[12740] = 12'b111111111111;
assign CPM[12741] = 12'b111111111111;
assign CPM[12742] = 12'b111111111111;
assign CPM[12743] = 12'b111111111111;
assign CPM[12744] = 12'b111111111111;
assign CPM[12745] = 12'b111111111111;
assign CPM[12746] = 12'b000000000000;
assign CPM[12747] = 12'b000000000000;
assign CPM[12748] = 12'b000000000000;
assign CPM[12749] = 12'b000000000000;
assign CPM[12750] = 12'b000000000000;
assign CPM[12751] = 12'b000000000000;
assign CPM[12752] = 12'b000000000000;
assign CPM[12753] = 12'b000000000000;
assign CPM[12754] = 12'b000000000000;
assign CPM[12755] = 12'b000000000000;
assign CPM[12756] = 12'b000000000000;
assign CPM[12757] = 12'b000000000000;
assign CPM[12758] = 12'b000000000000;
assign CPM[12759] = 12'b000000000000;
assign CPM[12760] = 12'b000000000000;
assign CPM[12761] = 12'b000000000000;
assign CPM[12762] = 12'b111111111111;
assign CPM[12763] = 12'b111111111111;
assign CPM[12764] = 12'b111111111111;
assign CPM[12765] = 12'b111111111111;
assign CPM[12766] = 12'b111111111111;
assign CPM[12767] = 12'b111111111111;
assign CPM[12768] = 12'b111111111111;
assign CPM[12769] = 12'b111111111111;
assign CPM[12770] = 12'b111111111111;
assign CPM[12771] = 12'b111111111111;
assign CPM[12772] = 12'b111111111111;
assign CPM[12773] = 12'b111111111111;
assign CPM[12774] = 12'b111111111111;
assign CPM[12775] = 12'b111111111111;
assign CPM[12776] = 12'b111111111111;
assign CPM[12777] = 12'b111111111111;
assign CPM[12778] = 12'b000000000000;
assign CPM[12779] = 12'b000000000000;
assign CPM[12780] = 12'b000000000000;
assign CPM[12781] = 12'b000000000000;
assign CPM[12782] = 12'b000000000000;
assign CPM[12783] = 12'b000000000000;
assign CPM[12784] = 12'b000000000000;
assign CPM[12785] = 12'b000000000000;
assign CPM[12786] = 12'b000000000000;
assign CPM[12787] = 12'b000000000000;
assign CPM[12788] = 12'b000000000000;
assign CPM[12789] = 12'b000000000000;
assign CPM[12790] = 12'b000000000000;
assign CPM[12791] = 12'b000000000000;
assign CPM[12792] = 12'b000000000000;
assign CPM[12793] = 12'b000000000000;
assign CPM[12794] = 12'b111111111111;
assign CPM[12795] = 12'b111111111111;
assign CPM[12796] = 12'b111111111111;
assign CPM[12797] = 12'b111111111111;
assign CPM[12798] = 12'b111111111111;
assign CPM[12799] = 12'b111111111111;
assign CPM[12800] = 12'b111111111111;
assign CPM[12801] = 12'b111111111111;
assign CPM[12802] = 12'b111111111111;
assign CPM[12803] = 12'b111111111111;
assign CPM[12804] = 12'b111111111111;
assign CPM[12805] = 12'b111111111111;
assign CPM[12806] = 12'b111111111111;
assign CPM[12807] = 12'b111111111111;
assign CPM[12808] = 12'b111111111111;
assign CPM[12809] = 12'b111111111111;
assign CPM[12810] = 12'b000000000000;
assign CPM[12811] = 12'b000000000000;
assign CPM[12812] = 12'b000000000000;
assign CPM[12813] = 12'b000000000000;
assign CPM[12814] = 12'b000000000000;
assign CPM[12815] = 12'b000000000000;
assign CPM[12816] = 12'b000000000000;
assign CPM[12817] = 12'b000000000000;
assign CPM[12818] = 12'b000000000000;
assign CPM[12819] = 12'b000000000000;
assign CPM[12820] = 12'b000000000000;
assign CPM[12821] = 12'b000000000000;
assign CPM[12822] = 12'b000000000000;
assign CPM[12823] = 12'b000000000000;
assign CPM[12824] = 12'b000000000000;
assign CPM[12825] = 12'b000000000000;
assign CPM[12826] = 12'b111111111111;
assign CPM[12827] = 12'b111111111111;
assign CPM[12828] = 12'b111111111111;
assign CPM[12829] = 12'b111111111111;
assign CPM[12830] = 12'b111111111111;
assign CPM[12831] = 12'b111111111111;
assign CPM[12832] = 12'b111111111111;
assign CPM[12833] = 12'b111111111111;
assign CPM[12834] = 12'b111111111111;
assign CPM[12835] = 12'b111111111111;
assign CPM[12836] = 12'b111111111111;
assign CPM[12837] = 12'b111111111111;
assign CPM[12838] = 12'b111111111111;
assign CPM[12839] = 12'b111111111111;
assign CPM[12840] = 12'b111111111111;
assign CPM[12841] = 12'b111111111111;
assign CPM[12842] = 12'b111111111111;
assign CPM[12843] = 12'b111111111111;
assign CPM[12844] = 12'b111111111111;
assign CPM[12845] = 12'b111111111111;
assign CPM[12846] = 12'b111111111111;
assign CPM[12847] = 12'b111111111111;
assign CPM[12848] = 12'b111111111111;
assign CPM[12849] = 12'b111111111111;
assign CPM[12850] = 12'b111111111111;
assign CPM[12851] = 12'b111111111111;
assign CPM[12852] = 12'b111111111111;
assign CPM[12853] = 12'b111111111111;
assign CPM[12854] = 12'b000000000000;
assign CPM[12855] = 12'b000000000000;
assign CPM[12856] = 12'b000000000000;
assign CPM[12857] = 12'b000000000000;
assign CPM[12858] = 12'b111111111111;
assign CPM[12859] = 12'b111111111111;
assign CPM[12860] = 12'b111111111111;
assign CPM[12861] = 12'b111111111111;
assign CPM[12862] = 12'b111111111111;
assign CPM[12863] = 12'b111111111111;
assign CPM[12864] = 12'b111111111111;
assign CPM[12865] = 12'b111111111111;
assign CPM[12866] = 12'b111111111111;
assign CPM[12867] = 12'b111111111111;
assign CPM[12868] = 12'b111111111111;
assign CPM[12869] = 12'b111111111111;
assign CPM[12870] = 12'b111111111111;
assign CPM[12871] = 12'b111111111111;
assign CPM[12872] = 12'b111111111111;
assign CPM[12873] = 12'b111111111111;
assign CPM[12874] = 12'b111111111111;
assign CPM[12875] = 12'b111111111111;
assign CPM[12876] = 12'b111111111111;
assign CPM[12877] = 12'b111111111111;
assign CPM[12878] = 12'b111111111111;
assign CPM[12879] = 12'b111111111111;
assign CPM[12880] = 12'b111111111111;
assign CPM[12881] = 12'b111111111111;
assign CPM[12882] = 12'b111111111111;
assign CPM[12883] = 12'b111111111111;
assign CPM[12884] = 12'b111111111111;
assign CPM[12885] = 12'b111111111111;
assign CPM[12886] = 12'b000000000000;
assign CPM[12887] = 12'b000000000000;
assign CPM[12888] = 12'b000000000000;
assign CPM[12889] = 12'b000000000000;
assign CPM[12890] = 12'b111111111111;
assign CPM[12891] = 12'b111111111111;
assign CPM[12892] = 12'b111111111111;
assign CPM[12893] = 12'b111111111111;
assign CPM[12894] = 12'b111111111111;
assign CPM[12895] = 12'b111111111111;
assign CPM[12896] = 12'b111111111111;
assign CPM[12897] = 12'b111111111111;
assign CPM[12898] = 12'b111111111111;
assign CPM[12899] = 12'b111111111111;
assign CPM[12900] = 12'b111111111111;
assign CPM[12901] = 12'b111111111111;
assign CPM[12902] = 12'b111111111111;
assign CPM[12903] = 12'b111111111111;
assign CPM[12904] = 12'b111111111111;
assign CPM[12905] = 12'b111111111111;
assign CPM[12906] = 12'b111111111111;
assign CPM[12907] = 12'b111111111111;
assign CPM[12908] = 12'b111111111111;
assign CPM[12909] = 12'b111111111111;
assign CPM[12910] = 12'b111111111111;
assign CPM[12911] = 12'b111111111111;
assign CPM[12912] = 12'b111111111111;
assign CPM[12913] = 12'b111111111111;
assign CPM[12914] = 12'b111111111111;
assign CPM[12915] = 12'b111111111111;
assign CPM[12916] = 12'b111111111111;
assign CPM[12917] = 12'b111111111111;
assign CPM[12918] = 12'b000000000000;
assign CPM[12919] = 12'b000000000000;
assign CPM[12920] = 12'b000000000000;
assign CPM[12921] = 12'b000000000000;
assign CPM[12922] = 12'b111111111111;
assign CPM[12923] = 12'b111111111111;
assign CPM[12924] = 12'b111111111111;
assign CPM[12925] = 12'b111111111111;
assign CPM[12926] = 12'b111111111111;
assign CPM[12927] = 12'b111111111111;
assign CPM[12928] = 12'b111111111111;
assign CPM[12929] = 12'b111111111111;
assign CPM[12930] = 12'b111111111111;
assign CPM[12931] = 12'b111111111111;
assign CPM[12932] = 12'b111111111111;
assign CPM[12933] = 12'b111111111111;
assign CPM[12934] = 12'b111111111111;
assign CPM[12935] = 12'b111111111111;
assign CPM[12936] = 12'b111111111111;
assign CPM[12937] = 12'b111111111111;
assign CPM[12938] = 12'b111111111111;
assign CPM[12939] = 12'b111111111111;
assign CPM[12940] = 12'b111111111111;
assign CPM[12941] = 12'b111111111111;
assign CPM[12942] = 12'b111111111111;
assign CPM[12943] = 12'b111111111111;
assign CPM[12944] = 12'b111111111111;
assign CPM[12945] = 12'b111111111111;
assign CPM[12946] = 12'b111111111111;
assign CPM[12947] = 12'b111111111111;
assign CPM[12948] = 12'b111111111111;
assign CPM[12949] = 12'b111111111111;
assign CPM[12950] = 12'b000000000000;
assign CPM[12951] = 12'b000000000000;
assign CPM[12952] = 12'b000000000000;
assign CPM[12953] = 12'b000000000000;
assign CPM[12954] = 12'b111111111111;
assign CPM[12955] = 12'b111111111111;
assign CPM[12956] = 12'b111111111111;
assign CPM[12957] = 12'b111111111111;
assign CPM[12958] = 12'b111111111111;
assign CPM[12959] = 12'b111111111111;
assign CPM[12960] = 12'b111111111111;
assign CPM[12961] = 12'b111111111111;
assign CPM[12962] = 12'b111111111111;
assign CPM[12963] = 12'b111111111111;
assign CPM[12964] = 12'b111111111111;
assign CPM[12965] = 12'b111111111111;
assign CPM[12966] = 12'b111111111111;
assign CPM[12967] = 12'b111111111111;
assign CPM[12968] = 12'b111111111111;
assign CPM[12969] = 12'b111111111111;
assign CPM[12970] = 12'b111111111111;
assign CPM[12971] = 12'b111111111111;
assign CPM[12972] = 12'b111111111111;
assign CPM[12973] = 12'b111111111111;
assign CPM[12974] = 12'b111111111111;
assign CPM[12975] = 12'b111111111111;
assign CPM[12976] = 12'b111111111111;
assign CPM[12977] = 12'b111111111111;
assign CPM[12978] = 12'b111111111111;
assign CPM[12979] = 12'b111111111111;
assign CPM[12980] = 12'b111111111111;
assign CPM[12981] = 12'b111111111111;
assign CPM[12982] = 12'b000000000000;
assign CPM[12983] = 12'b000000000000;
assign CPM[12984] = 12'b000000000000;
assign CPM[12985] = 12'b000000000000;
assign CPM[12986] = 12'b111111111111;
assign CPM[12987] = 12'b111111111111;
assign CPM[12988] = 12'b111111111111;
assign CPM[12989] = 12'b111111111111;
assign CPM[12990] = 12'b111111111111;
assign CPM[12991] = 12'b111111111111;
assign CPM[12992] = 12'b111111111111;
assign CPM[12993] = 12'b111111111111;
assign CPM[12994] = 12'b111111111111;
assign CPM[12995] = 12'b111111111111;
assign CPM[12996] = 12'b111111111111;
assign CPM[12997] = 12'b111111111111;
assign CPM[12998] = 12'b000000000000;
assign CPM[12999] = 12'b000000000000;
assign CPM[13000] = 12'b000000000000;
assign CPM[13001] = 12'b000000000000;
assign CPM[13002] = 12'b111111111111;
assign CPM[13003] = 12'b111111111111;
assign CPM[13004] = 12'b111111111111;
assign CPM[13005] = 12'b111111111111;
assign CPM[13006] = 12'b111111111111;
assign CPM[13007] = 12'b111111111111;
assign CPM[13008] = 12'b111111111111;
assign CPM[13009] = 12'b111111111111;
assign CPM[13010] = 12'b111111111111;
assign CPM[13011] = 12'b111111111111;
assign CPM[13012] = 12'b111111111111;
assign CPM[13013] = 12'b111111111111;
assign CPM[13014] = 12'b000000000000;
assign CPM[13015] = 12'b000000000000;
assign CPM[13016] = 12'b000000000000;
assign CPM[13017] = 12'b000000000000;
assign CPM[13018] = 12'b111111111111;
assign CPM[13019] = 12'b111111111111;
assign CPM[13020] = 12'b111111111111;
assign CPM[13021] = 12'b111111111111;
assign CPM[13022] = 12'b111111111111;
assign CPM[13023] = 12'b111111111111;
assign CPM[13024] = 12'b111111111111;
assign CPM[13025] = 12'b111111111111;
assign CPM[13026] = 12'b111111111111;
assign CPM[13027] = 12'b111111111111;
assign CPM[13028] = 12'b111111111111;
assign CPM[13029] = 12'b111111111111;
assign CPM[13030] = 12'b000000000000;
assign CPM[13031] = 12'b000000000000;
assign CPM[13032] = 12'b000000000000;
assign CPM[13033] = 12'b000000000000;
assign CPM[13034] = 12'b111111111111;
assign CPM[13035] = 12'b111111111111;
assign CPM[13036] = 12'b111111111111;
assign CPM[13037] = 12'b111111111111;
assign CPM[13038] = 12'b111111111111;
assign CPM[13039] = 12'b111111111111;
assign CPM[13040] = 12'b111111111111;
assign CPM[13041] = 12'b111111111111;
assign CPM[13042] = 12'b111111111111;
assign CPM[13043] = 12'b111111111111;
assign CPM[13044] = 12'b111111111111;
assign CPM[13045] = 12'b111111111111;
assign CPM[13046] = 12'b000000000000;
assign CPM[13047] = 12'b000000000000;
assign CPM[13048] = 12'b000000000000;
assign CPM[13049] = 12'b000000000000;
assign CPM[13050] = 12'b111111111111;
assign CPM[13051] = 12'b111111111111;
assign CPM[13052] = 12'b111111111111;
assign CPM[13053] = 12'b111111111111;
assign CPM[13054] = 12'b111111111111;
assign CPM[13055] = 12'b111111111111;
assign CPM[13056] = 12'b111111111111;
assign CPM[13057] = 12'b111111111111;
assign CPM[13058] = 12'b111111111111;
assign CPM[13059] = 12'b111111111111;
assign CPM[13060] = 12'b111111111111;
assign CPM[13061] = 12'b111111111111;
assign CPM[13062] = 12'b000000000000;
assign CPM[13063] = 12'b000000000000;
assign CPM[13064] = 12'b000000000000;
assign CPM[13065] = 12'b000000000000;
assign CPM[13066] = 12'b111111111111;
assign CPM[13067] = 12'b111111111111;
assign CPM[13068] = 12'b111111111111;
assign CPM[13069] = 12'b111111111111;
assign CPM[13070] = 12'b111111111111;
assign CPM[13071] = 12'b111111111111;
assign CPM[13072] = 12'b111111111111;
assign CPM[13073] = 12'b111111111111;
assign CPM[13074] = 12'b111111111111;
assign CPM[13075] = 12'b111111111111;
assign CPM[13076] = 12'b111111111111;
assign CPM[13077] = 12'b111111111111;
assign CPM[13078] = 12'b000000000000;
assign CPM[13079] = 12'b000000000000;
assign CPM[13080] = 12'b000000000000;
assign CPM[13081] = 12'b000000000000;
assign CPM[13082] = 12'b111111111111;
assign CPM[13083] = 12'b111111111111;
assign CPM[13084] = 12'b111111111111;
assign CPM[13085] = 12'b111111111111;
assign CPM[13086] = 12'b111111111111;
assign CPM[13087] = 12'b111111111111;
assign CPM[13088] = 12'b111111111111;
assign CPM[13089] = 12'b111111111111;
assign CPM[13090] = 12'b111111111111;
assign CPM[13091] = 12'b111111111111;
assign CPM[13092] = 12'b111111111111;
assign CPM[13093] = 12'b111111111111;
assign CPM[13094] = 12'b000000000000;
assign CPM[13095] = 12'b000000000000;
assign CPM[13096] = 12'b000000000000;
assign CPM[13097] = 12'b000000000000;
assign CPM[13098] = 12'b111111111111;
assign CPM[13099] = 12'b111111111111;
assign CPM[13100] = 12'b111111111111;
assign CPM[13101] = 12'b111111111111;
assign CPM[13102] = 12'b111111111111;
assign CPM[13103] = 12'b111111111111;
assign CPM[13104] = 12'b111111111111;
assign CPM[13105] = 12'b111111111111;
assign CPM[13106] = 12'b111111111111;
assign CPM[13107] = 12'b111111111111;
assign CPM[13108] = 12'b111111111111;
assign CPM[13109] = 12'b111111111111;
assign CPM[13110] = 12'b000000000000;
assign CPM[13111] = 12'b000000000000;
assign CPM[13112] = 12'b000000000000;
assign CPM[13113] = 12'b000000000000;
assign CPM[13114] = 12'b111111111111;
assign CPM[13115] = 12'b111111111111;
assign CPM[13116] = 12'b111111111111;
assign CPM[13117] = 12'b111111111111;
assign CPM[13118] = 12'b111111111111;
assign CPM[13119] = 12'b111111111111;
assign CPM[13120] = 12'b111111111111;
assign CPM[13121] = 12'b111111111111;
assign CPM[13122] = 12'b111111111111;
assign CPM[13123] = 12'b111111111111;
assign CPM[13124] = 12'b111111111111;
assign CPM[13125] = 12'b111111111111;
assign CPM[13126] = 12'b111111111111;
assign CPM[13127] = 12'b111111111111;
assign CPM[13128] = 12'b111111111111;
assign CPM[13129] = 12'b111111111111;
assign CPM[13130] = 12'b000000000000;
assign CPM[13131] = 12'b000000000000;
assign CPM[13132] = 12'b000000000000;
assign CPM[13133] = 12'b000000000000;
assign CPM[13134] = 12'b000000000000;
assign CPM[13135] = 12'b000000000000;
assign CPM[13136] = 12'b000000000000;
assign CPM[13137] = 12'b000000000000;
assign CPM[13138] = 12'b000000000000;
assign CPM[13139] = 12'b000000000000;
assign CPM[13140] = 12'b000000000000;
assign CPM[13141] = 12'b000000000000;
assign CPM[13142] = 12'b111111111111;
assign CPM[13143] = 12'b111111111111;
assign CPM[13144] = 12'b111111111111;
assign CPM[13145] = 12'b111111111111;
assign CPM[13146] = 12'b111111111111;
assign CPM[13147] = 12'b111111111111;
assign CPM[13148] = 12'b111111111111;
assign CPM[13149] = 12'b111111111111;
assign CPM[13150] = 12'b111111111111;
assign CPM[13151] = 12'b111111111111;
assign CPM[13152] = 12'b111111111111;
assign CPM[13153] = 12'b111111111111;
assign CPM[13154] = 12'b111111111111;
assign CPM[13155] = 12'b111111111111;
assign CPM[13156] = 12'b111111111111;
assign CPM[13157] = 12'b111111111111;
assign CPM[13158] = 12'b111111111111;
assign CPM[13159] = 12'b111111111111;
assign CPM[13160] = 12'b111111111111;
assign CPM[13161] = 12'b111111111111;
assign CPM[13162] = 12'b000000000000;
assign CPM[13163] = 12'b000000000000;
assign CPM[13164] = 12'b000000000000;
assign CPM[13165] = 12'b000000000000;
assign CPM[13166] = 12'b000000000000;
assign CPM[13167] = 12'b000000000000;
assign CPM[13168] = 12'b000000000000;
assign CPM[13169] = 12'b000000000000;
assign CPM[13170] = 12'b000000000000;
assign CPM[13171] = 12'b000000000000;
assign CPM[13172] = 12'b000000000000;
assign CPM[13173] = 12'b000000000000;
assign CPM[13174] = 12'b111111111111;
assign CPM[13175] = 12'b111111111111;
assign CPM[13176] = 12'b111111111111;
assign CPM[13177] = 12'b111111111111;
assign CPM[13178] = 12'b111111111111;
assign CPM[13179] = 12'b111111111111;
assign CPM[13180] = 12'b111111111111;
assign CPM[13181] = 12'b111111111111;
assign CPM[13182] = 12'b111111111111;
assign CPM[13183] = 12'b111111111111;
assign CPM[13184] = 12'b111111111111;
assign CPM[13185] = 12'b111111111111;
assign CPM[13186] = 12'b111111111111;
assign CPM[13187] = 12'b111111111111;
assign CPM[13188] = 12'b111111111111;
assign CPM[13189] = 12'b111111111111;
assign CPM[13190] = 12'b111111111111;
assign CPM[13191] = 12'b111111111111;
assign CPM[13192] = 12'b111111111111;
assign CPM[13193] = 12'b111111111111;
assign CPM[13194] = 12'b000000000000;
assign CPM[13195] = 12'b000000000000;
assign CPM[13196] = 12'b000000000000;
assign CPM[13197] = 12'b000000000000;
assign CPM[13198] = 12'b000000000000;
assign CPM[13199] = 12'b000000000000;
assign CPM[13200] = 12'b000000000000;
assign CPM[13201] = 12'b000000000000;
assign CPM[13202] = 12'b000000000000;
assign CPM[13203] = 12'b000000000000;
assign CPM[13204] = 12'b000000000000;
assign CPM[13205] = 12'b000000000000;
assign CPM[13206] = 12'b111111111111;
assign CPM[13207] = 12'b111111111111;
assign CPM[13208] = 12'b111111111111;
assign CPM[13209] = 12'b111111111111;
assign CPM[13210] = 12'b111111111111;
assign CPM[13211] = 12'b111111111111;
assign CPM[13212] = 12'b111111111111;
assign CPM[13213] = 12'b111111111111;
assign CPM[13214] = 12'b111111111111;
assign CPM[13215] = 12'b111111111111;
assign CPM[13216] = 12'b111111111111;
assign CPM[13217] = 12'b111111111111;
assign CPM[13218] = 12'b111111111111;
assign CPM[13219] = 12'b111111111111;
assign CPM[13220] = 12'b111111111111;
assign CPM[13221] = 12'b111111111111;
assign CPM[13222] = 12'b111111111111;
assign CPM[13223] = 12'b111111111111;
assign CPM[13224] = 12'b111111111111;
assign CPM[13225] = 12'b111111111111;
assign CPM[13226] = 12'b000000000000;
assign CPM[13227] = 12'b000000000000;
assign CPM[13228] = 12'b000000000000;
assign CPM[13229] = 12'b000000000000;
assign CPM[13230] = 12'b000000000000;
assign CPM[13231] = 12'b000000000000;
assign CPM[13232] = 12'b000000000000;
assign CPM[13233] = 12'b000000000000;
assign CPM[13234] = 12'b000000000000;
assign CPM[13235] = 12'b000000000000;
assign CPM[13236] = 12'b000000000000;
assign CPM[13237] = 12'b000000000000;
assign CPM[13238] = 12'b111111111111;
assign CPM[13239] = 12'b111111111111;
assign CPM[13240] = 12'b111111111111;
assign CPM[13241] = 12'b111111111111;
assign CPM[13242] = 12'b111111111111;
assign CPM[13243] = 12'b111111111111;
assign CPM[13244] = 12'b111111111111;
assign CPM[13245] = 12'b111111111111;
assign CPM[13246] = 12'b111111111111;
assign CPM[13247] = 12'b111111111111;
assign CPM[13248] = 12'b111111111111;
assign CPM[13249] = 12'b111111111111;
assign CPM[13250] = 12'b111111111111;
assign CPM[13251] = 12'b111111111111;
assign CPM[13252] = 12'b111111111111;
assign CPM[13253] = 12'b111111111111;
assign CPM[13254] = 12'b111111111111;
assign CPM[13255] = 12'b111111111111;
assign CPM[13256] = 12'b111111111111;
assign CPM[13257] = 12'b111111111111;
assign CPM[13258] = 12'b111111111111;
assign CPM[13259] = 12'b111111111111;
assign CPM[13260] = 12'b111111111111;
assign CPM[13261] = 12'b111111111111;
assign CPM[13262] = 12'b111111111111;
assign CPM[13263] = 12'b111111111111;
assign CPM[13264] = 12'b111111111111;
assign CPM[13265] = 12'b111111111111;
assign CPM[13266] = 12'b111111111111;
assign CPM[13267] = 12'b111111111111;
assign CPM[13268] = 12'b111111111111;
assign CPM[13269] = 12'b111111111111;
assign CPM[13270] = 12'b111111111111;
assign CPM[13271] = 12'b111111111111;
assign CPM[13272] = 12'b111111111111;
assign CPM[13273] = 12'b111111111111;
assign CPM[13274] = 12'b111111111111;
assign CPM[13275] = 12'b111111111111;
assign CPM[13276] = 12'b111111111111;
assign CPM[13277] = 12'b111111111111;
assign CPM[13278] = 12'b111111111111;
assign CPM[13279] = 12'b111111111111;
assign CPM[13280] = 12'b111111111111;
assign CPM[13281] = 12'b111111111111;
assign CPM[13282] = 12'b111111111111;
assign CPM[13283] = 12'b111111111111;
assign CPM[13284] = 12'b111111111111;
assign CPM[13285] = 12'b111111111111;
assign CPM[13286] = 12'b111111111111;
assign CPM[13287] = 12'b111111111111;
assign CPM[13288] = 12'b111111111111;
assign CPM[13289] = 12'b111111111111;
assign CPM[13290] = 12'b111111111111;
assign CPM[13291] = 12'b111111111111;
assign CPM[13292] = 12'b111111111111;
assign CPM[13293] = 12'b111111111111;
assign CPM[13294] = 12'b111111111111;
assign CPM[13295] = 12'b111111111111;
assign CPM[13296] = 12'b111111111111;
assign CPM[13297] = 12'b111111111111;
assign CPM[13298] = 12'b111111111111;
assign CPM[13299] = 12'b111111111111;
assign CPM[13300] = 12'b111111111111;
assign CPM[13301] = 12'b111111111111;
assign CPM[13302] = 12'b111111111111;
assign CPM[13303] = 12'b111111111111;
assign CPM[13304] = 12'b111111111111;
assign CPM[13305] = 12'b111111111111;
assign CPM[13306] = 12'b111111111111;
assign CPM[13307] = 12'b111111111111;
assign CPM[13308] = 12'b111111111111;
assign CPM[13309] = 12'b111111111111;
assign CPM[13310] = 12'b111111111111;
assign CPM[13311] = 12'b111111111111;

endmodule
