`timescale 1ns/1ps

module q3_t();

    reg clk = 0;
    reg rst_n = 0;
    wire [8-1:0] out;

    parameter cyc = 10;
    always #(cyc/2) clk = ~clk;

    Q4 M1(
        .clk(clk),
        .rst_n(rst_n),
        .out(out)
    );

    initial begin
        $dumpfile("q3.vcd");
        $dumpvars("+all");
    end
    initial begin
        @(negedge clk)
        rst_n = 1;
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        @(negedge clk)
        $finish;
    end



endmodule
