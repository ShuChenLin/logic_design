`timescale 1ns/1ps

module fpga1(clk, 
