`timescale 1ns/1ps

module mem_addr_gen(
   input clk,
   input rst,
   input [9:0] h_cnt,
   input [9:0] v_cnt,
   input [8:0] word_num,
   input [5:0] letter,
   input correct,
   input [10:0] word_cnt,
   output reg [3:0] red, green, blue
   );
    
   wire [11:0] Upperletter [1663:0];
   wire [11:0] Lowerletter [1663:0];
   wire [11:0] otherletter [255:0];
   wire [15:0] place, place2, place3;
   
   assign place = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * letter);
   assign place2 = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * (letter - 26));
   assign place3 = (h_cnt % 8) + 8*(v_cnt % 8) + (64 * (letter - 30));
   
   always @(*) begin
        {red, green, blue} = 12'b111111111111;
        if (h_cnt >= 80 && h_cnt <= 560 && v_cnt >= 208 && v_cnt <= 280) begin
            if (word_num > 298 || (v_cnt / 8) == 27 || (v_cnt) / 8 == 29 || (v_cnt) / 8 == 31 || (v_cnt) / 8 == 33 || (v_cnt) / 8 == 35) {red, green, blue} = 12'b111111111111;
            else begin
                if (correct && word_num == word_cnt) begin
                    if (letter <= 25) {red, green, blue} = (Lowerletter[place] == 12'b111111111111) ? 12'b111111111111 : 12'b111100000000;
                    else if (letter >= 26 && letter <= 29) {red, green, blue} = (otherletter[place2] == 12'b111111111111) ? 12'b111111111111 : 12'b111100000000;
                    else {red, green, blue} = (Upperletter[place3] == 12'b111111111111) ? 12'b111111111111 : 12'b111100000000;
                end else if (word_num < word_cnt) begin
                    if (letter <= 25) {red, green, blue} = (Lowerletter[place] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;
                    else if (letter >= 26 && letter <= 29) {red, green, blue} = (otherletter[place2] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;
                    else {red, green, blue} = (Upperletter[place3] == 12'b111111111111) ? 12'b111111111111 : 12'b000011110000;
                end else begin
                    if (letter <= 25) {red, green, blue} = Lowerletter[place];
                    else if (letter >= 26 && letter <= 29) {red, green, blue} = otherletter[place2];
                    else {red, green, blue} = Upperletter[place3];
                end
            end
//            {red, green, blue} = Upperletter[0];
        end
    end
    
assign otherletter[0] = 12'b111111111111;
assign otherletter[1] = 12'b111111111111;
assign otherletter[2] = 12'b111111111111;
assign otherletter[3] = 12'b111111111111;
assign otherletter[4] = 12'b111111111111;
assign otherletter[5] = 12'b111111111111;
assign otherletter[6] = 12'b111111111111;
assign otherletter[7] = 12'b111111111111;
assign otherletter[8] = 12'b111111111111;
assign otherletter[9] = 12'b111111111111;
assign otherletter[10] = 12'b111111111111;
assign otherletter[11] = 12'b111111111111;
assign otherletter[12] = 12'b111111111111;
assign otherletter[13] = 12'b111111111111;
assign otherletter[14] = 12'b111111111111;
assign otherletter[15] = 12'b111111111111;
assign otherletter[16] = 12'b111111111111;
assign otherletter[17] = 12'b111111111111;
assign otherletter[18] = 12'b111111111111;
assign otherletter[19] = 12'b111111111111;
assign otherletter[20] = 12'b111111111111;
assign otherletter[21] = 12'b111111111111;
assign otherletter[22] = 12'b111111111111;
assign otherletter[23] = 12'b111111111111;
assign otherletter[24] = 12'b111111111111;
assign otherletter[25] = 12'b111111111111;
assign otherletter[26] = 12'b111111111111;
assign otherletter[27] = 12'b111111111111;
assign otherletter[28] = 12'b111111111111;
assign otherletter[29] = 12'b111111111111;
assign otherletter[30] = 12'b111111111111;
assign otherletter[31] = 12'b111111111111;
assign otherletter[32] = 12'b111111111111;
assign otherletter[33] = 12'b111111111111;
assign otherletter[34] = 12'b111111111111;
assign otherletter[35] = 12'b111111111111;
assign otherletter[36] = 12'b111111111111;
assign otherletter[37] = 12'b111111111111;
assign otherletter[38] = 12'b111111111111;
assign otherletter[39] = 12'b111111111111;
assign otherletter[40] = 12'b111111111111;
assign otherletter[41] = 12'b111111111111;
assign otherletter[42] = 12'b111111111111;
assign otherletter[43] = 12'b111111111111;
assign otherletter[44] = 12'b111111111111;
assign otherletter[45] = 12'b111111111111;
assign otherletter[46] = 12'b111111111111;
assign otherletter[47] = 12'b111111111111;
assign otherletter[48] = 12'b111111111111;
assign otherletter[49] = 12'b111111111111;
assign otherletter[50] = 12'b111111111111;
assign otherletter[51] = 12'b111111111111;
assign otherletter[52] = 12'b111111111111;
assign otherletter[53] = 12'b111111111111;
assign otherletter[54] = 12'b111111111111;
assign otherletter[55] = 12'b111111111111;
assign otherletter[56] = 12'b111111111111;
assign otherletter[57] = 12'b111111111111;
assign otherletter[58] = 12'b111111111111;
assign otherletter[59] = 12'b111111111111;
assign otherletter[60] = 12'b111111111111;
assign otherletter[61] = 12'b111111111111;
assign otherletter[62] = 12'b111111111111;
assign otherletter[63] = 12'b111111111111;
assign otherletter[64] = 12'b111111111111;
assign otherletter[65] = 12'b111111111111;
assign otherletter[66] = 12'b111111111111;
assign otherletter[67] = 12'b111111111111;
assign otherletter[68] = 12'b111111111111;
assign otherletter[69] = 12'b111111111111;
assign otherletter[70] = 12'b111111111111;
assign otherletter[71] = 12'b111111111111;
assign otherletter[72] = 12'b111111111111;
assign otherletter[73] = 12'b111111111111;
assign otherletter[74] = 12'b111111111111;
assign otherletter[75] = 12'b111111111111;
assign otherletter[76] = 12'b111111111111;
assign otherletter[77] = 12'b111111111111;
assign otherletter[78] = 12'b111111111111;
assign otherletter[79] = 12'b111111111111;
assign otherletter[80] = 12'b111111111111;
assign otherletter[81] = 12'b111111111111;
assign otherletter[82] = 12'b111111111111;
assign otherletter[83] = 12'b111111111111;
assign otherletter[84] = 12'b111111111111;
assign otherletter[85] = 12'b111111111111;
assign otherletter[86] = 12'b111111111111;
assign otherletter[87] = 12'b111111111111;
assign otherletter[88] = 12'b111111111111;
assign otherletter[89] = 12'b111111111111;
assign otherletter[90] = 12'b111111111111;
assign otherletter[91] = 12'b111111111111;
assign otherletter[92] = 12'b111111111111;
assign otherletter[93] = 12'b111111111111;
assign otherletter[94] = 12'b111111111111;
assign otherletter[95] = 12'b111111111111;
assign otherletter[96] = 12'b111111111111;
assign otherletter[97] = 12'b111111111111;
assign otherletter[98] = 12'b111111111111;
assign otherletter[99] = 12'b111111111111;
assign otherletter[100] = 12'b111111111111;
assign otherletter[101] = 12'b111111111111;
assign otherletter[102] = 12'b111111111111;
assign otherletter[103] = 12'b111111111111;
assign otherletter[104] = 12'b111111111111;
assign otherletter[105] = 12'b111111111111;
assign otherletter[106] = 12'b111111111111;
assign otherletter[107] = 12'b111111111111;
assign otherletter[108] = 12'b111111111111;
assign otherletter[109] = 12'b111111111111;
assign otherletter[110] = 12'b111111111111;
assign otherletter[111] = 12'b111111111111;
assign otherletter[112] = 12'b111111111111;
assign otherletter[113] = 12'b111111111111;
assign otherletter[114] = 12'b111111111111;
assign otherletter[115] = 12'b000000000000;
assign otherletter[116] = 12'b111111111111;
assign otherletter[117] = 12'b111111111111;
assign otherletter[118] = 12'b111111111111;
assign otherletter[119] = 12'b111111111111;
assign otherletter[120] = 12'b111111111111;
assign otherletter[121] = 12'b111111111111;
assign otherletter[122] = 12'b111111111111;
assign otherletter[123] = 12'b000000000000;
assign otherletter[124] = 12'b111111111111;
assign otherletter[125] = 12'b111111111111;
assign otherletter[126] = 12'b111111111111;
assign otherletter[127] = 12'b111111111111;
assign otherletter[128] = 12'b111111111111;
assign otherletter[129] = 12'b111111111111;
assign otherletter[130] = 12'b111111111111;
assign otherletter[131] = 12'b111111111111;
assign otherletter[132] = 12'b111111111111;
assign otherletter[133] = 12'b111111111111;
assign otherletter[134] = 12'b111111111111;
assign otherletter[135] = 12'b111111111111;
assign otherletter[136] = 12'b111111111111;
assign otherletter[137] = 12'b111111111111;
assign otherletter[138] = 12'b111111111111;
assign otherletter[139] = 12'b111111111111;
assign otherletter[140] = 12'b111111111111;
assign otherletter[141] = 12'b111111111111;
assign otherletter[142] = 12'b111111111111;
assign otherletter[143] = 12'b111111111111;
assign otherletter[144] = 12'b111111111111;
assign otherletter[145] = 12'b111111111111;
assign otherletter[146] = 12'b111111111111;
assign otherletter[147] = 12'b111111111111;
assign otherletter[148] = 12'b111111111111;
assign otherletter[149] = 12'b111111111111;
assign otherletter[150] = 12'b111111111111;
assign otherletter[151] = 12'b111111111111;
assign otherletter[152] = 12'b111111111111;
assign otherletter[153] = 12'b111111111111;
assign otherletter[154] = 12'b111111111111;
assign otherletter[155] = 12'b111111111111;
assign otherletter[156] = 12'b111111111111;
assign otherletter[157] = 12'b111111111111;
assign otherletter[158] = 12'b111111111111;
assign otherletter[159] = 12'b111111111111;
assign otherletter[160] = 12'b111111111111;
assign otherletter[161] = 12'b111111111111;
assign otherletter[162] = 12'b111111111111;
assign otherletter[163] = 12'b111111111111;
assign otherletter[164] = 12'b111111111111;
assign otherletter[165] = 12'b111111111111;
assign otherletter[166] = 12'b111111111111;
assign otherletter[167] = 12'b111111111111;
assign otherletter[168] = 12'b111111111111;
assign otherletter[169] = 12'b111111111111;
assign otherletter[170] = 12'b111111111111;
assign otherletter[171] = 12'b111111111111;
assign otherletter[172] = 12'b111111111111;
assign otherletter[173] = 12'b111111111111;
assign otherletter[174] = 12'b111111111111;
assign otherletter[175] = 12'b111111111111;
assign otherletter[176] = 12'b111111111111;
assign otherletter[177] = 12'b111111111111;
assign otherletter[178] = 12'b111111111111;
assign otherletter[179] = 12'b000000000000;
assign otherletter[180] = 12'b111111111111;
assign otherletter[181] = 12'b111111111111;
assign otherletter[182] = 12'b111111111111;
assign otherletter[183] = 12'b111111111111;
assign otherletter[184] = 12'b111111111111;
assign otherletter[185] = 12'b111111111111;
assign otherletter[186] = 12'b111111111111;
assign otherletter[187] = 12'b111111111111;
assign otherletter[188] = 12'b111111111111;
assign otherletter[189] = 12'b111111111111;
assign otherletter[190] = 12'b111111111111;
assign otherletter[191] = 12'b111111111111;
assign otherletter[192] = 12'b111111111111;
assign otherletter[193] = 12'b111111111111;
assign otherletter[194] = 12'b111111111111;
assign otherletter[195] = 12'b000000000000;
assign otherletter[196] = 12'b111111111111;
assign otherletter[197] = 12'b111111111111;
assign otherletter[198] = 12'b111111111111;
assign otherletter[199] = 12'b111111111111;
assign otherletter[200] = 12'b111111111111;
assign otherletter[201] = 12'b111111111111;
assign otherletter[202] = 12'b111111111111;
assign otherletter[203] = 12'b000000000000;
assign otherletter[204] = 12'b111111111111;
assign otherletter[205] = 12'b111111111111;
assign otherletter[206] = 12'b111111111111;
assign otherletter[207] = 12'b111111111111;
assign otherletter[208] = 12'b111111111111;
assign otherletter[209] = 12'b111111111111;
assign otherletter[210] = 12'b111111111111;
assign otherletter[211] = 12'b111111111111;
assign otherletter[212] = 12'b111111111111;
assign otherletter[213] = 12'b111111111111;
assign otherletter[214] = 12'b111111111111;
assign otherletter[215] = 12'b111111111111;
assign otherletter[216] = 12'b111111111111;
assign otherletter[217] = 12'b111111111111;
assign otherletter[218] = 12'b111111111111;
assign otherletter[219] = 12'b111111111111;
assign otherletter[220] = 12'b111111111111;
assign otherletter[221] = 12'b111111111111;
assign otherletter[222] = 12'b111111111111;
assign otherletter[223] = 12'b111111111111;
assign otherletter[224] = 12'b111111111111;
assign otherletter[225] = 12'b111111111111;
assign otherletter[226] = 12'b111111111111;
assign otherletter[227] = 12'b111111111111;
assign otherletter[228] = 12'b111111111111;
assign otherletter[229] = 12'b111111111111;
assign otherletter[230] = 12'b111111111111;
assign otherletter[231] = 12'b111111111111;
assign otherletter[232] = 12'b111111111111;
assign otherletter[233] = 12'b111111111111;
assign otherletter[234] = 12'b111111111111;
assign otherletter[235] = 12'b111111111111;
assign otherletter[236] = 12'b111111111111;
assign otherletter[237] = 12'b111111111111;
assign otherletter[238] = 12'b111111111111;
assign otherletter[239] = 12'b111111111111;
assign otherletter[240] = 12'b111111111111;
assign otherletter[241] = 12'b111111111111;
assign otherletter[242] = 12'b111111111111;
assign otherletter[243] = 12'b111111111111;
assign otherletter[244] = 12'b111111111111;
assign otherletter[245] = 12'b111111111111;
assign otherletter[246] = 12'b111111111111;
assign otherletter[247] = 12'b111111111111;
assign otherletter[248] = 12'b111111111111;
assign otherletter[249] = 12'b111111111111;
assign otherletter[250] = 12'b111111111111;
assign otherletter[251] = 12'b111111111111;
assign otherletter[252] = 12'b111111111111;
assign otherletter[253] = 12'b111111111111;
assign otherletter[254] = 12'b111111111111;
assign otherletter[255] = 12'b111111111111;    
assign Lowerletter[0] = 12'b111111111111;
assign Lowerletter[1] = 12'b111111111111;
assign Lowerletter[2] = 12'b111111111111;
assign Lowerletter[3] = 12'b111111111111;
assign Lowerletter[4] = 12'b111111111111;
assign Lowerletter[5] = 12'b111111111111;
assign Lowerletter[6] = 12'b111111111111;
assign Lowerletter[7] = 12'b111111111111;
assign Lowerletter[8] = 12'b111111111111;
assign Lowerletter[9] = 12'b111111111111;
assign Lowerletter[10] = 12'b111111111111;
assign Lowerletter[11] = 12'b111111111111;
assign Lowerletter[12] = 12'b111111111111;
assign Lowerletter[13] = 12'b111111111111;
assign Lowerletter[14] = 12'b111111111111;
assign Lowerletter[15] = 12'b111111111111;
assign Lowerletter[16] = 12'b111111111111;
assign Lowerletter[17] = 12'b111111111111;
assign Lowerletter[18] = 12'b000000000000;
assign Lowerletter[19] = 12'b000000000000;
assign Lowerletter[20] = 12'b000000000000;
assign Lowerletter[21] = 12'b111111111111;
assign Lowerletter[22] = 12'b111111111111;
assign Lowerletter[23] = 12'b111111111111;
assign Lowerletter[24] = 12'b111111111111;
assign Lowerletter[25] = 12'b111111111111;
assign Lowerletter[26] = 12'b111111111111;
assign Lowerletter[27] = 12'b111111111111;
assign Lowerletter[28] = 12'b111111111111;
assign Lowerletter[29] = 12'b000000000000;
assign Lowerletter[30] = 12'b111111111111;
assign Lowerletter[31] = 12'b111111111111;
assign Lowerletter[32] = 12'b111111111111;
assign Lowerletter[33] = 12'b111111111111;
assign Lowerletter[34] = 12'b111111111111;
assign Lowerletter[35] = 12'b000000000000;
assign Lowerletter[36] = 12'b000000000000;
assign Lowerletter[37] = 12'b000000000000;
assign Lowerletter[38] = 12'b111111111111;
assign Lowerletter[39] = 12'b111111111111;
assign Lowerletter[40] = 12'b111111111111;
assign Lowerletter[41] = 12'b111111111111;
assign Lowerletter[42] = 12'b000000000000;
assign Lowerletter[43] = 12'b111111111111;
assign Lowerletter[44] = 12'b111111111111;
assign Lowerletter[45] = 12'b000000000000;
assign Lowerletter[46] = 12'b111111111111;
assign Lowerletter[47] = 12'b111111111111;
assign Lowerletter[48] = 12'b111111111111;
assign Lowerletter[49] = 12'b111111111111;
assign Lowerletter[50] = 12'b111111111111;
assign Lowerletter[51] = 12'b000000000000;
assign Lowerletter[52] = 12'b000000000000;
assign Lowerletter[53] = 12'b000000000000;
assign Lowerletter[54] = 12'b111111111111;
assign Lowerletter[55] = 12'b111111111111;
assign Lowerletter[56] = 12'b111111111111;
assign Lowerletter[57] = 12'b111111111111;
assign Lowerletter[58] = 12'b111111111111;
assign Lowerletter[59] = 12'b111111111111;
assign Lowerletter[60] = 12'b111111111111;
assign Lowerletter[61] = 12'b111111111111;
assign Lowerletter[62] = 12'b111111111111;
assign Lowerletter[63] = 12'b111111111111;
assign Lowerletter[64] = 12'b111111111111;
assign Lowerletter[65] = 12'b111111111111;
assign Lowerletter[66] = 12'b000000000000;
assign Lowerletter[67] = 12'b111111111111;
assign Lowerletter[68] = 12'b111111111111;
assign Lowerletter[69] = 12'b111111111111;
assign Lowerletter[70] = 12'b111111111111;
assign Lowerletter[71] = 12'b111111111111;
assign Lowerletter[72] = 12'b111111111111;
assign Lowerletter[73] = 12'b111111111111;
assign Lowerletter[74] = 12'b000000000000;
assign Lowerletter[75] = 12'b111111111111;
assign Lowerletter[76] = 12'b111111111111;
assign Lowerletter[77] = 12'b111111111111;
assign Lowerletter[78] = 12'b111111111111;
assign Lowerletter[79] = 12'b111111111111;
assign Lowerletter[80] = 12'b111111111111;
assign Lowerletter[81] = 12'b111111111111;
assign Lowerletter[82] = 12'b000000000000;
assign Lowerletter[83] = 12'b111111111111;
assign Lowerletter[84] = 12'b111111111111;
assign Lowerletter[85] = 12'b111111111111;
assign Lowerletter[86] = 12'b111111111111;
assign Lowerletter[87] = 12'b111111111111;
assign Lowerletter[88] = 12'b111111111111;
assign Lowerletter[89] = 12'b111111111111;
assign Lowerletter[90] = 12'b000000000000;
assign Lowerletter[91] = 12'b111111111111;
assign Lowerletter[92] = 12'b000000000000;
assign Lowerletter[93] = 12'b111111111111;
assign Lowerletter[94] = 12'b111111111111;
assign Lowerletter[95] = 12'b111111111111;
assign Lowerletter[96] = 12'b111111111111;
assign Lowerletter[97] = 12'b111111111111;
assign Lowerletter[98] = 12'b000000000000;
assign Lowerletter[99] = 12'b000000000000;
assign Lowerletter[100] = 12'b111111111111;
assign Lowerletter[101] = 12'b000000000000;
assign Lowerletter[102] = 12'b111111111111;
assign Lowerletter[103] = 12'b111111111111;
assign Lowerletter[104] = 12'b111111111111;
assign Lowerletter[105] = 12'b111111111111;
assign Lowerletter[106] = 12'b000000000000;
assign Lowerletter[107] = 12'b111111111111;
assign Lowerletter[108] = 12'b111111111111;
assign Lowerletter[109] = 12'b000000000000;
assign Lowerletter[110] = 12'b111111111111;
assign Lowerletter[111] = 12'b111111111111;
assign Lowerletter[112] = 12'b111111111111;
assign Lowerletter[113] = 12'b111111111111;
assign Lowerletter[114] = 12'b000000000000;
assign Lowerletter[115] = 12'b000000000000;
assign Lowerletter[116] = 12'b000000000000;
assign Lowerletter[117] = 12'b111111111111;
assign Lowerletter[118] = 12'b111111111111;
assign Lowerletter[119] = 12'b111111111111;
assign Lowerletter[120] = 12'b111111111111;
assign Lowerletter[121] = 12'b111111111111;
assign Lowerletter[122] = 12'b111111111111;
assign Lowerletter[123] = 12'b111111111111;
assign Lowerletter[124] = 12'b111111111111;
assign Lowerletter[125] = 12'b111111111111;
assign Lowerletter[126] = 12'b111111111111;
assign Lowerletter[127] = 12'b111111111111;
assign Lowerletter[128] = 12'b111111111111;
assign Lowerletter[129] = 12'b111111111111;
assign Lowerletter[130] = 12'b111111111111;
assign Lowerletter[131] = 12'b111111111111;
assign Lowerletter[132] = 12'b111111111111;
assign Lowerletter[133] = 12'b111111111111;
assign Lowerletter[134] = 12'b111111111111;
assign Lowerletter[135] = 12'b111111111111;
assign Lowerletter[136] = 12'b111111111111;
assign Lowerletter[137] = 12'b111111111111;
assign Lowerletter[138] = 12'b111111111111;
assign Lowerletter[139] = 12'b111111111111;
assign Lowerletter[140] = 12'b111111111111;
assign Lowerletter[141] = 12'b111111111111;
assign Lowerletter[142] = 12'b111111111111;
assign Lowerletter[143] = 12'b111111111111;
assign Lowerletter[144] = 12'b111111111111;
assign Lowerletter[145] = 12'b111111111111;
assign Lowerletter[146] = 12'b111111111111;
assign Lowerletter[147] = 12'b000000000000;
assign Lowerletter[148] = 12'b000000000000;
assign Lowerletter[149] = 12'b111111111111;
assign Lowerletter[150] = 12'b111111111111;
assign Lowerletter[151] = 12'b111111111111;
assign Lowerletter[152] = 12'b111111111111;
assign Lowerletter[153] = 12'b111111111111;
assign Lowerletter[154] = 12'b000000000000;
assign Lowerletter[155] = 12'b111111111111;
assign Lowerletter[156] = 12'b111111111111;
assign Lowerletter[157] = 12'b000000000000;
assign Lowerletter[158] = 12'b111111111111;
assign Lowerletter[159] = 12'b111111111111;
assign Lowerletter[160] = 12'b111111111111;
assign Lowerletter[161] = 12'b111111111111;
assign Lowerletter[162] = 12'b000000000000;
assign Lowerletter[163] = 12'b111111111111;
assign Lowerletter[164] = 12'b111111111111;
assign Lowerletter[165] = 12'b111111111111;
assign Lowerletter[166] = 12'b111111111111;
assign Lowerletter[167] = 12'b111111111111;
assign Lowerletter[168] = 12'b111111111111;
assign Lowerletter[169] = 12'b111111111111;
assign Lowerletter[170] = 12'b000000000000;
assign Lowerletter[171] = 12'b111111111111;
assign Lowerletter[172] = 12'b111111111111;
assign Lowerletter[173] = 12'b000000000000;
assign Lowerletter[174] = 12'b111111111111;
assign Lowerletter[175] = 12'b111111111111;
assign Lowerletter[176] = 12'b111111111111;
assign Lowerletter[177] = 12'b111111111111;
assign Lowerletter[178] = 12'b111111111111;
assign Lowerletter[179] = 12'b000000000000;
assign Lowerletter[180] = 12'b000000000000;
assign Lowerletter[181] = 12'b111111111111;
assign Lowerletter[182] = 12'b111111111111;
assign Lowerletter[183] = 12'b111111111111;
assign Lowerletter[184] = 12'b111111111111;
assign Lowerletter[185] = 12'b111111111111;
assign Lowerletter[186] = 12'b111111111111;
assign Lowerletter[187] = 12'b111111111111;
assign Lowerletter[188] = 12'b111111111111;
assign Lowerletter[189] = 12'b111111111111;
assign Lowerletter[190] = 12'b111111111111;
assign Lowerletter[191] = 12'b111111111111;
assign Lowerletter[192] = 12'b111111111111;
assign Lowerletter[193] = 12'b111111111111;
assign Lowerletter[194] = 12'b111111111111;
assign Lowerletter[195] = 12'b111111111111;
assign Lowerletter[196] = 12'b111111111111;
assign Lowerletter[197] = 12'b000000000000;
assign Lowerletter[198] = 12'b111111111111;
assign Lowerletter[199] = 12'b111111111111;
assign Lowerletter[200] = 12'b111111111111;
assign Lowerletter[201] = 12'b111111111111;
assign Lowerletter[202] = 12'b111111111111;
assign Lowerletter[203] = 12'b111111111111;
assign Lowerletter[204] = 12'b111111111111;
assign Lowerletter[205] = 12'b000000000000;
assign Lowerletter[206] = 12'b111111111111;
assign Lowerletter[207] = 12'b111111111111;
assign Lowerletter[208] = 12'b111111111111;
assign Lowerletter[209] = 12'b111111111111;
assign Lowerletter[210] = 12'b111111111111;
assign Lowerletter[211] = 12'b111111111111;
assign Lowerletter[212] = 12'b111111111111;
assign Lowerletter[213] = 12'b000000000000;
assign Lowerletter[214] = 12'b111111111111;
assign Lowerletter[215] = 12'b111111111111;
assign Lowerletter[216] = 12'b111111111111;
assign Lowerletter[217] = 12'b111111111111;
assign Lowerletter[218] = 12'b111111111111;
assign Lowerletter[219] = 12'b000000000000;
assign Lowerletter[220] = 12'b000000000000;
assign Lowerletter[221] = 12'b000000000000;
assign Lowerletter[222] = 12'b111111111111;
assign Lowerletter[223] = 12'b111111111111;
assign Lowerletter[224] = 12'b111111111111;
assign Lowerletter[225] = 12'b111111111111;
assign Lowerletter[226] = 12'b000000000000;
assign Lowerletter[227] = 12'b111111111111;
assign Lowerletter[228] = 12'b111111111111;
assign Lowerletter[229] = 12'b000000000000;
assign Lowerletter[230] = 12'b111111111111;
assign Lowerletter[231] = 12'b111111111111;
assign Lowerletter[232] = 12'b111111111111;
assign Lowerletter[233] = 12'b111111111111;
assign Lowerletter[234] = 12'b000000000000;
assign Lowerletter[235] = 12'b111111111111;
assign Lowerletter[236] = 12'b111111111111;
assign Lowerletter[237] = 12'b000000000000;
assign Lowerletter[238] = 12'b111111111111;
assign Lowerletter[239] = 12'b111111111111;
assign Lowerletter[240] = 12'b111111111111;
assign Lowerletter[241] = 12'b111111111111;
assign Lowerletter[242] = 12'b000000000000;
assign Lowerletter[243] = 12'b000000000000;
assign Lowerletter[244] = 12'b000000000000;
assign Lowerletter[245] = 12'b000000000000;
assign Lowerletter[246] = 12'b111111111111;
assign Lowerletter[247] = 12'b111111111111;
assign Lowerletter[248] = 12'b111111111111;
assign Lowerletter[249] = 12'b111111111111;
assign Lowerletter[250] = 12'b111111111111;
assign Lowerletter[251] = 12'b111111111111;
assign Lowerletter[252] = 12'b111111111111;
assign Lowerletter[253] = 12'b111111111111;
assign Lowerletter[254] = 12'b111111111111;
assign Lowerletter[255] = 12'b111111111111;
assign Lowerletter[256] = 12'b111111111111;
assign Lowerletter[257] = 12'b111111111111;
assign Lowerletter[258] = 12'b111111111111;
assign Lowerletter[259] = 12'b111111111111;
assign Lowerletter[260] = 12'b111111111111;
assign Lowerletter[261] = 12'b111111111111;
assign Lowerletter[262] = 12'b111111111111;
assign Lowerletter[263] = 12'b111111111111;
assign Lowerletter[264] = 12'b111111111111;
assign Lowerletter[265] = 12'b111111111111;
assign Lowerletter[266] = 12'b111111111111;
assign Lowerletter[267] = 12'b111111111111;
assign Lowerletter[268] = 12'b111111111111;
assign Lowerletter[269] = 12'b111111111111;
assign Lowerletter[270] = 12'b111111111111;
assign Lowerletter[271] = 12'b111111111111;
assign Lowerletter[272] = 12'b111111111111;
assign Lowerletter[273] = 12'b111111111111;
assign Lowerletter[274] = 12'b111111111111;
assign Lowerletter[275] = 12'b000000000000;
assign Lowerletter[276] = 12'b000000000000;
assign Lowerletter[277] = 12'b000000000000;
assign Lowerletter[278] = 12'b111111111111;
assign Lowerletter[279] = 12'b111111111111;
assign Lowerletter[280] = 12'b111111111111;
assign Lowerletter[281] = 12'b111111111111;
assign Lowerletter[282] = 12'b000000000000;
assign Lowerletter[283] = 12'b111111111111;
assign Lowerletter[284] = 12'b111111111111;
assign Lowerletter[285] = 12'b000000000000;
assign Lowerletter[286] = 12'b111111111111;
assign Lowerletter[287] = 12'b111111111111;
assign Lowerletter[288] = 12'b111111111111;
assign Lowerletter[289] = 12'b111111111111;
assign Lowerletter[290] = 12'b000000000000;
assign Lowerletter[291] = 12'b000000000000;
assign Lowerletter[292] = 12'b000000000000;
assign Lowerletter[293] = 12'b111111111111;
assign Lowerletter[294] = 12'b111111111111;
assign Lowerletter[295] = 12'b111111111111;
assign Lowerletter[296] = 12'b111111111111;
assign Lowerletter[297] = 12'b111111111111;
assign Lowerletter[298] = 12'b000000000000;
assign Lowerletter[299] = 12'b111111111111;
assign Lowerletter[300] = 12'b111111111111;
assign Lowerletter[301] = 12'b111111111111;
assign Lowerletter[302] = 12'b111111111111;
assign Lowerletter[303] = 12'b111111111111;
assign Lowerletter[304] = 12'b111111111111;
assign Lowerletter[305] = 12'b111111111111;
assign Lowerletter[306] = 12'b111111111111;
assign Lowerletter[307] = 12'b000000000000;
assign Lowerletter[308] = 12'b000000000000;
assign Lowerletter[309] = 12'b000000000000;
assign Lowerletter[310] = 12'b111111111111;
assign Lowerletter[311] = 12'b111111111111;
assign Lowerletter[312] = 12'b111111111111;
assign Lowerletter[313] = 12'b111111111111;
assign Lowerletter[314] = 12'b111111111111;
assign Lowerletter[315] = 12'b111111111111;
assign Lowerletter[316] = 12'b111111111111;
assign Lowerletter[317] = 12'b111111111111;
assign Lowerletter[318] = 12'b111111111111;
assign Lowerletter[319] = 12'b111111111111;
assign Lowerletter[320] = 12'b111111111111;
assign Lowerletter[321] = 12'b111111111111;
assign Lowerletter[322] = 12'b111111111111;
assign Lowerletter[323] = 12'b000000000000;
assign Lowerletter[324] = 12'b000000000000;
assign Lowerletter[325] = 12'b111111111111;
assign Lowerletter[326] = 12'b111111111111;
assign Lowerletter[327] = 12'b111111111111;
assign Lowerletter[328] = 12'b111111111111;
assign Lowerletter[329] = 12'b111111111111;
assign Lowerletter[330] = 12'b111111111111;
assign Lowerletter[331] = 12'b000000000000;
assign Lowerletter[332] = 12'b111111111111;
assign Lowerletter[333] = 12'b111111111111;
assign Lowerletter[334] = 12'b111111111111;
assign Lowerletter[335] = 12'b111111111111;
assign Lowerletter[336] = 12'b111111111111;
assign Lowerletter[337] = 12'b111111111111;
assign Lowerletter[338] = 12'b000000000000;
assign Lowerletter[339] = 12'b000000000000;
assign Lowerletter[340] = 12'b000000000000;
assign Lowerletter[341] = 12'b000000000000;
assign Lowerletter[342] = 12'b111111111111;
assign Lowerletter[343] = 12'b111111111111;
assign Lowerletter[344] = 12'b111111111111;
assign Lowerletter[345] = 12'b111111111111;
assign Lowerletter[346] = 12'b111111111111;
assign Lowerletter[347] = 12'b000000000000;
assign Lowerletter[348] = 12'b111111111111;
assign Lowerletter[349] = 12'b111111111111;
assign Lowerletter[350] = 12'b111111111111;
assign Lowerletter[351] = 12'b111111111111;
assign Lowerletter[352] = 12'b111111111111;
assign Lowerletter[353] = 12'b111111111111;
assign Lowerletter[354] = 12'b111111111111;
assign Lowerletter[355] = 12'b000000000000;
assign Lowerletter[356] = 12'b111111111111;
assign Lowerletter[357] = 12'b111111111111;
assign Lowerletter[358] = 12'b111111111111;
assign Lowerletter[359] = 12'b111111111111;
assign Lowerletter[360] = 12'b111111111111;
assign Lowerletter[361] = 12'b111111111111;
assign Lowerletter[362] = 12'b111111111111;
assign Lowerletter[363] = 12'b000000000000;
assign Lowerletter[364] = 12'b111111111111;
assign Lowerletter[365] = 12'b111111111111;
assign Lowerletter[366] = 12'b111111111111;
assign Lowerletter[367] = 12'b111111111111;
assign Lowerletter[368] = 12'b111111111111;
assign Lowerletter[369] = 12'b111111111111;
assign Lowerletter[370] = 12'b111111111111;
assign Lowerletter[371] = 12'b000000000000;
assign Lowerletter[372] = 12'b111111111111;
assign Lowerletter[373] = 12'b111111111111;
assign Lowerletter[374] = 12'b111111111111;
assign Lowerletter[375] = 12'b111111111111;
assign Lowerletter[376] = 12'b111111111111;
assign Lowerletter[377] = 12'b111111111111;
assign Lowerletter[378] = 12'b111111111111;
assign Lowerletter[379] = 12'b111111111111;
assign Lowerletter[380] = 12'b111111111111;
assign Lowerletter[381] = 12'b111111111111;
assign Lowerletter[382] = 12'b111111111111;
assign Lowerletter[383] = 12'b111111111111;
assign Lowerletter[384] = 12'b111111111111;
assign Lowerletter[385] = 12'b111111111111;
assign Lowerletter[386] = 12'b111111111111;
assign Lowerletter[387] = 12'b111111111111;
assign Lowerletter[388] = 12'b111111111111;
assign Lowerletter[389] = 12'b111111111111;
assign Lowerletter[390] = 12'b111111111111;
assign Lowerletter[391] = 12'b111111111111;
assign Lowerletter[392] = 12'b111111111111;
assign Lowerletter[393] = 12'b111111111111;
assign Lowerletter[394] = 12'b111111111111;
assign Lowerletter[395] = 12'b111111111111;
assign Lowerletter[396] = 12'b111111111111;
assign Lowerletter[397] = 12'b111111111111;
assign Lowerletter[398] = 12'b111111111111;
assign Lowerletter[399] = 12'b111111111111;
assign Lowerletter[400] = 12'b111111111111;
assign Lowerletter[401] = 12'b111111111111;
assign Lowerletter[402] = 12'b111111111111;
assign Lowerletter[403] = 12'b000000000000;
assign Lowerletter[404] = 12'b000000000000;
assign Lowerletter[405] = 12'b000000000000;
assign Lowerletter[406] = 12'b111111111111;
assign Lowerletter[407] = 12'b111111111111;
assign Lowerletter[408] = 12'b111111111111;
assign Lowerletter[409] = 12'b111111111111;
assign Lowerletter[410] = 12'b000000000000;
assign Lowerletter[411] = 12'b111111111111;
assign Lowerletter[412] = 12'b111111111111;
assign Lowerletter[413] = 12'b000000000000;
assign Lowerletter[414] = 12'b111111111111;
assign Lowerletter[415] = 12'b111111111111;
assign Lowerletter[416] = 12'b111111111111;
assign Lowerletter[417] = 12'b111111111111;
assign Lowerletter[418] = 12'b111111111111;
assign Lowerletter[419] = 12'b000000000000;
assign Lowerletter[420] = 12'b000000000000;
assign Lowerletter[421] = 12'b000000000000;
assign Lowerletter[422] = 12'b111111111111;
assign Lowerletter[423] = 12'b111111111111;
assign Lowerletter[424] = 12'b111111111111;
assign Lowerletter[425] = 12'b111111111111;
assign Lowerletter[426] = 12'b111111111111;
assign Lowerletter[427] = 12'b111111111111;
assign Lowerletter[428] = 12'b111111111111;
assign Lowerletter[429] = 12'b000000000000;
assign Lowerletter[430] = 12'b111111111111;
assign Lowerletter[431] = 12'b111111111111;
assign Lowerletter[432] = 12'b111111111111;
assign Lowerletter[433] = 12'b111111111111;
assign Lowerletter[434] = 12'b000000000000;
assign Lowerletter[435] = 12'b111111111111;
assign Lowerletter[436] = 12'b111111111111;
assign Lowerletter[437] = 12'b000000000000;
assign Lowerletter[438] = 12'b111111111111;
assign Lowerletter[439] = 12'b111111111111;
assign Lowerletter[440] = 12'b111111111111;
assign Lowerletter[441] = 12'b111111111111;
assign Lowerletter[442] = 12'b111111111111;
assign Lowerletter[443] = 12'b000000000000;
assign Lowerletter[444] = 12'b000000000000;
assign Lowerletter[445] = 12'b111111111111;
assign Lowerletter[446] = 12'b111111111111;
assign Lowerletter[447] = 12'b111111111111;
assign Lowerletter[448] = 12'b111111111111;
assign Lowerletter[449] = 12'b111111111111;
assign Lowerletter[450] = 12'b000000000000;
assign Lowerletter[451] = 12'b111111111111;
assign Lowerletter[452] = 12'b111111111111;
assign Lowerletter[453] = 12'b111111111111;
assign Lowerletter[454] = 12'b111111111111;
assign Lowerletter[455] = 12'b111111111111;
assign Lowerletter[456] = 12'b111111111111;
assign Lowerletter[457] = 12'b111111111111;
assign Lowerletter[458] = 12'b000000000000;
assign Lowerletter[459] = 12'b111111111111;
assign Lowerletter[460] = 12'b111111111111;
assign Lowerletter[461] = 12'b111111111111;
assign Lowerletter[462] = 12'b111111111111;
assign Lowerletter[463] = 12'b111111111111;
assign Lowerletter[464] = 12'b111111111111;
assign Lowerletter[465] = 12'b111111111111;
assign Lowerletter[466] = 12'b000000000000;
assign Lowerletter[467] = 12'b111111111111;
assign Lowerletter[468] = 12'b111111111111;
assign Lowerletter[469] = 12'b111111111111;
assign Lowerletter[470] = 12'b111111111111;
assign Lowerletter[471] = 12'b111111111111;
assign Lowerletter[472] = 12'b111111111111;
assign Lowerletter[473] = 12'b111111111111;
assign Lowerletter[474] = 12'b000000000000;
assign Lowerletter[475] = 12'b111111111111;
assign Lowerletter[476] = 12'b000000000000;
assign Lowerletter[477] = 12'b111111111111;
assign Lowerletter[478] = 12'b111111111111;
assign Lowerletter[479] = 12'b111111111111;
assign Lowerletter[480] = 12'b111111111111;
assign Lowerletter[481] = 12'b111111111111;
assign Lowerletter[482] = 12'b000000000000;
assign Lowerletter[483] = 12'b000000000000;
assign Lowerletter[484] = 12'b111111111111;
assign Lowerletter[485] = 12'b000000000000;
assign Lowerletter[486] = 12'b111111111111;
assign Lowerletter[487] = 12'b111111111111;
assign Lowerletter[488] = 12'b111111111111;
assign Lowerletter[489] = 12'b111111111111;
assign Lowerletter[490] = 12'b000000000000;
assign Lowerletter[491] = 12'b111111111111;
assign Lowerletter[492] = 12'b111111111111;
assign Lowerletter[493] = 12'b000000000000;
assign Lowerletter[494] = 12'b111111111111;
assign Lowerletter[495] = 12'b111111111111;
assign Lowerletter[496] = 12'b111111111111;
assign Lowerletter[497] = 12'b111111111111;
assign Lowerletter[498] = 12'b000000000000;
assign Lowerletter[499] = 12'b111111111111;
assign Lowerletter[500] = 12'b111111111111;
assign Lowerletter[501] = 12'b000000000000;
assign Lowerletter[502] = 12'b111111111111;
assign Lowerletter[503] = 12'b111111111111;
assign Lowerletter[504] = 12'b111111111111;
assign Lowerletter[505] = 12'b111111111111;
assign Lowerletter[506] = 12'b111111111111;
assign Lowerletter[507] = 12'b111111111111;
assign Lowerletter[508] = 12'b111111111111;
assign Lowerletter[509] = 12'b111111111111;
assign Lowerletter[510] = 12'b111111111111;
assign Lowerletter[511] = 12'b111111111111;
assign Lowerletter[512] = 12'b111111111111;
assign Lowerletter[513] = 12'b111111111111;
assign Lowerletter[514] = 12'b111111111111;
assign Lowerletter[515] = 12'b111111111111;
assign Lowerletter[516] = 12'b111111111111;
assign Lowerletter[517] = 12'b111111111111;
assign Lowerletter[518] = 12'b111111111111;
assign Lowerletter[519] = 12'b111111111111;
assign Lowerletter[520] = 12'b111111111111;
assign Lowerletter[521] = 12'b111111111111;
assign Lowerletter[522] = 12'b111111111111;
assign Lowerletter[523] = 12'b000000000000;
assign Lowerletter[524] = 12'b111111111111;
assign Lowerletter[525] = 12'b111111111111;
assign Lowerletter[526] = 12'b111111111111;
assign Lowerletter[527] = 12'b111111111111;
assign Lowerletter[528] = 12'b111111111111;
assign Lowerletter[529] = 12'b111111111111;
assign Lowerletter[530] = 12'b111111111111;
assign Lowerletter[531] = 12'b111111111111;
assign Lowerletter[532] = 12'b111111111111;
assign Lowerletter[533] = 12'b111111111111;
assign Lowerletter[534] = 12'b111111111111;
assign Lowerletter[535] = 12'b111111111111;
assign Lowerletter[536] = 12'b111111111111;
assign Lowerletter[537] = 12'b111111111111;
assign Lowerletter[538] = 12'b111111111111;
assign Lowerletter[539] = 12'b000000000000;
assign Lowerletter[540] = 12'b111111111111;
assign Lowerletter[541] = 12'b111111111111;
assign Lowerletter[542] = 12'b111111111111;
assign Lowerletter[543] = 12'b111111111111;
assign Lowerletter[544] = 12'b111111111111;
assign Lowerletter[545] = 12'b111111111111;
assign Lowerletter[546] = 12'b111111111111;
assign Lowerletter[547] = 12'b000000000000;
assign Lowerletter[548] = 12'b111111111111;
assign Lowerletter[549] = 12'b111111111111;
assign Lowerletter[550] = 12'b111111111111;
assign Lowerletter[551] = 12'b111111111111;
assign Lowerletter[552] = 12'b111111111111;
assign Lowerletter[553] = 12'b111111111111;
assign Lowerletter[554] = 12'b111111111111;
assign Lowerletter[555] = 12'b000000000000;
assign Lowerletter[556] = 12'b111111111111;
assign Lowerletter[557] = 12'b111111111111;
assign Lowerletter[558] = 12'b111111111111;
assign Lowerletter[559] = 12'b111111111111;
assign Lowerletter[560] = 12'b111111111111;
assign Lowerletter[561] = 12'b111111111111;
assign Lowerletter[562] = 12'b111111111111;
assign Lowerletter[563] = 12'b000000000000;
assign Lowerletter[564] = 12'b111111111111;
assign Lowerletter[565] = 12'b111111111111;
assign Lowerletter[566] = 12'b111111111111;
assign Lowerletter[567] = 12'b111111111111;
assign Lowerletter[568] = 12'b111111111111;
assign Lowerletter[569] = 12'b111111111111;
assign Lowerletter[570] = 12'b111111111111;
assign Lowerletter[571] = 12'b111111111111;
assign Lowerletter[572] = 12'b111111111111;
assign Lowerletter[573] = 12'b111111111111;
assign Lowerletter[574] = 12'b111111111111;
assign Lowerletter[575] = 12'b111111111111;
assign Lowerletter[576] = 12'b111111111111;
assign Lowerletter[577] = 12'b111111111111;
assign Lowerletter[578] = 12'b111111111111;
assign Lowerletter[579] = 12'b111111111111;
assign Lowerletter[580] = 12'b111111111111;
assign Lowerletter[581] = 12'b111111111111;
assign Lowerletter[582] = 12'b111111111111;
assign Lowerletter[583] = 12'b111111111111;
assign Lowerletter[584] = 12'b111111111111;
assign Lowerletter[585] = 12'b111111111111;
assign Lowerletter[586] = 12'b111111111111;
assign Lowerletter[587] = 12'b111111111111;
assign Lowerletter[588] = 12'b111111111111;
assign Lowerletter[589] = 12'b111111111111;
assign Lowerletter[590] = 12'b111111111111;
assign Lowerletter[591] = 12'b111111111111;
assign Lowerletter[592] = 12'b111111111111;
assign Lowerletter[593] = 12'b111111111111;
assign Lowerletter[594] = 12'b111111111111;
assign Lowerletter[595] = 12'b111111111111;
assign Lowerletter[596] = 12'b000000000000;
assign Lowerletter[597] = 12'b111111111111;
assign Lowerletter[598] = 12'b111111111111;
assign Lowerletter[599] = 12'b111111111111;
assign Lowerletter[600] = 12'b111111111111;
assign Lowerletter[601] = 12'b111111111111;
assign Lowerletter[602] = 12'b111111111111;
assign Lowerletter[603] = 12'b111111111111;
assign Lowerletter[604] = 12'b111111111111;
assign Lowerletter[605] = 12'b111111111111;
assign Lowerletter[606] = 12'b111111111111;
assign Lowerletter[607] = 12'b111111111111;
assign Lowerletter[608] = 12'b111111111111;
assign Lowerletter[609] = 12'b111111111111;
assign Lowerletter[610] = 12'b111111111111;
assign Lowerletter[611] = 12'b111111111111;
assign Lowerletter[612] = 12'b000000000000;
assign Lowerletter[613] = 12'b111111111111;
assign Lowerletter[614] = 12'b111111111111;
assign Lowerletter[615] = 12'b111111111111;
assign Lowerletter[616] = 12'b111111111111;
assign Lowerletter[617] = 12'b111111111111;
assign Lowerletter[618] = 12'b111111111111;
assign Lowerletter[619] = 12'b111111111111;
assign Lowerletter[620] = 12'b000000000000;
assign Lowerletter[621] = 12'b111111111111;
assign Lowerletter[622] = 12'b111111111111;
assign Lowerletter[623] = 12'b111111111111;
assign Lowerletter[624] = 12'b111111111111;
assign Lowerletter[625] = 12'b111111111111;
assign Lowerletter[626] = 12'b000000000000;
assign Lowerletter[627] = 12'b111111111111;
assign Lowerletter[628] = 12'b000000000000;
assign Lowerletter[629] = 12'b111111111111;
assign Lowerletter[630] = 12'b111111111111;
assign Lowerletter[631] = 12'b111111111111;
assign Lowerletter[632] = 12'b111111111111;
assign Lowerletter[633] = 12'b111111111111;
assign Lowerletter[634] = 12'b111111111111;
assign Lowerletter[635] = 12'b000000000000;
assign Lowerletter[636] = 12'b111111111111;
assign Lowerletter[637] = 12'b111111111111;
assign Lowerletter[638] = 12'b111111111111;
assign Lowerletter[639] = 12'b111111111111;
assign Lowerletter[640] = 12'b111111111111;
assign Lowerletter[641] = 12'b111111111111;
assign Lowerletter[642] = 12'b000000000000;
assign Lowerletter[643] = 12'b111111111111;
assign Lowerletter[644] = 12'b111111111111;
assign Lowerletter[645] = 12'b111111111111;
assign Lowerletter[646] = 12'b111111111111;
assign Lowerletter[647] = 12'b111111111111;
assign Lowerletter[648] = 12'b111111111111;
assign Lowerletter[649] = 12'b111111111111;
assign Lowerletter[650] = 12'b000000000000;
assign Lowerletter[651] = 12'b111111111111;
assign Lowerletter[652] = 12'b111111111111;
assign Lowerletter[653] = 12'b111111111111;
assign Lowerletter[654] = 12'b111111111111;
assign Lowerletter[655] = 12'b111111111111;
assign Lowerletter[656] = 12'b111111111111;
assign Lowerletter[657] = 12'b111111111111;
assign Lowerletter[658] = 12'b000000000000;
assign Lowerletter[659] = 12'b111111111111;
assign Lowerletter[660] = 12'b111111111111;
assign Lowerletter[661] = 12'b000000000000;
assign Lowerletter[662] = 12'b111111111111;
assign Lowerletter[663] = 12'b111111111111;
assign Lowerletter[664] = 12'b111111111111;
assign Lowerletter[665] = 12'b111111111111;
assign Lowerletter[666] = 12'b000000000000;
assign Lowerletter[667] = 12'b111111111111;
assign Lowerletter[668] = 12'b000000000000;
assign Lowerletter[669] = 12'b111111111111;
assign Lowerletter[670] = 12'b111111111111;
assign Lowerletter[671] = 12'b111111111111;
assign Lowerletter[672] = 12'b111111111111;
assign Lowerletter[673] = 12'b111111111111;
assign Lowerletter[674] = 12'b000000000000;
assign Lowerletter[675] = 12'b000000000000;
assign Lowerletter[676] = 12'b111111111111;
assign Lowerletter[677] = 12'b111111111111;
assign Lowerletter[678] = 12'b111111111111;
assign Lowerletter[679] = 12'b111111111111;
assign Lowerletter[680] = 12'b111111111111;
assign Lowerletter[681] = 12'b111111111111;
assign Lowerletter[682] = 12'b000000000000;
assign Lowerletter[683] = 12'b111111111111;
assign Lowerletter[684] = 12'b000000000000;
assign Lowerletter[685] = 12'b111111111111;
assign Lowerletter[686] = 12'b111111111111;
assign Lowerletter[687] = 12'b111111111111;
assign Lowerletter[688] = 12'b111111111111;
assign Lowerletter[689] = 12'b111111111111;
assign Lowerletter[690] = 12'b000000000000;
assign Lowerletter[691] = 12'b111111111111;
assign Lowerletter[692] = 12'b111111111111;
assign Lowerletter[693] = 12'b000000000000;
assign Lowerletter[694] = 12'b111111111111;
assign Lowerletter[695] = 12'b111111111111;
assign Lowerletter[696] = 12'b111111111111;
assign Lowerletter[697] = 12'b111111111111;
assign Lowerletter[698] = 12'b111111111111;
assign Lowerletter[699] = 12'b111111111111;
assign Lowerletter[700] = 12'b111111111111;
assign Lowerletter[701] = 12'b111111111111;
assign Lowerletter[702] = 12'b111111111111;
assign Lowerletter[703] = 12'b111111111111;
assign Lowerletter[704] = 12'b111111111111;
assign Lowerletter[705] = 12'b111111111111;
assign Lowerletter[706] = 12'b111111111111;
assign Lowerletter[707] = 12'b000000000000;
assign Lowerletter[708] = 12'b111111111111;
assign Lowerletter[709] = 12'b111111111111;
assign Lowerletter[710] = 12'b111111111111;
assign Lowerletter[711] = 12'b111111111111;
assign Lowerletter[712] = 12'b111111111111;
assign Lowerletter[713] = 12'b111111111111;
assign Lowerletter[714] = 12'b111111111111;
assign Lowerletter[715] = 12'b000000000000;
assign Lowerletter[716] = 12'b111111111111;
assign Lowerletter[717] = 12'b111111111111;
assign Lowerletter[718] = 12'b111111111111;
assign Lowerletter[719] = 12'b111111111111;
assign Lowerletter[720] = 12'b111111111111;
assign Lowerletter[721] = 12'b111111111111;
assign Lowerletter[722] = 12'b111111111111;
assign Lowerletter[723] = 12'b000000000000;
assign Lowerletter[724] = 12'b111111111111;
assign Lowerletter[725] = 12'b111111111111;
assign Lowerletter[726] = 12'b111111111111;
assign Lowerletter[727] = 12'b111111111111;
assign Lowerletter[728] = 12'b111111111111;
assign Lowerletter[729] = 12'b111111111111;
assign Lowerletter[730] = 12'b111111111111;
assign Lowerletter[731] = 12'b000000000000;
assign Lowerletter[732] = 12'b111111111111;
assign Lowerletter[733] = 12'b111111111111;
assign Lowerletter[734] = 12'b111111111111;
assign Lowerletter[735] = 12'b111111111111;
assign Lowerletter[736] = 12'b111111111111;
assign Lowerletter[737] = 12'b111111111111;
assign Lowerletter[738] = 12'b111111111111;
assign Lowerletter[739] = 12'b000000000000;
assign Lowerletter[740] = 12'b111111111111;
assign Lowerletter[741] = 12'b111111111111;
assign Lowerletter[742] = 12'b111111111111;
assign Lowerletter[743] = 12'b111111111111;
assign Lowerletter[744] = 12'b111111111111;
assign Lowerletter[745] = 12'b111111111111;
assign Lowerletter[746] = 12'b111111111111;
assign Lowerletter[747] = 12'b000000000000;
assign Lowerletter[748] = 12'b111111111111;
assign Lowerletter[749] = 12'b111111111111;
assign Lowerletter[750] = 12'b111111111111;
assign Lowerletter[751] = 12'b111111111111;
assign Lowerletter[752] = 12'b111111111111;
assign Lowerletter[753] = 12'b111111111111;
assign Lowerletter[754] = 12'b111111111111;
assign Lowerletter[755] = 12'b000000000000;
assign Lowerletter[756] = 12'b111111111111;
assign Lowerletter[757] = 12'b111111111111;
assign Lowerletter[758] = 12'b111111111111;
assign Lowerletter[759] = 12'b111111111111;
assign Lowerletter[760] = 12'b111111111111;
assign Lowerletter[761] = 12'b111111111111;
assign Lowerletter[762] = 12'b111111111111;
assign Lowerletter[763] = 12'b111111111111;
assign Lowerletter[764] = 12'b111111111111;
assign Lowerletter[765] = 12'b111111111111;
assign Lowerletter[766] = 12'b111111111111;
assign Lowerletter[767] = 12'b111111111111;
assign Lowerletter[768] = 12'b111111111111;
assign Lowerletter[769] = 12'b111111111111;
assign Lowerletter[770] = 12'b111111111111;
assign Lowerletter[771] = 12'b111111111111;
assign Lowerletter[772] = 12'b111111111111;
assign Lowerletter[773] = 12'b111111111111;
assign Lowerletter[774] = 12'b111111111111;
assign Lowerletter[775] = 12'b111111111111;
assign Lowerletter[776] = 12'b111111111111;
assign Lowerletter[777] = 12'b111111111111;
assign Lowerletter[778] = 12'b111111111111;
assign Lowerletter[779] = 12'b111111111111;
assign Lowerletter[780] = 12'b111111111111;
assign Lowerletter[781] = 12'b111111111111;
assign Lowerletter[782] = 12'b111111111111;
assign Lowerletter[783] = 12'b111111111111;
assign Lowerletter[784] = 12'b111111111111;
assign Lowerletter[785] = 12'b000000000000;
assign Lowerletter[786] = 12'b000000000000;
assign Lowerletter[787] = 12'b111111111111;
assign Lowerletter[788] = 12'b000000000000;
assign Lowerletter[789] = 12'b111111111111;
assign Lowerletter[790] = 12'b111111111111;
assign Lowerletter[791] = 12'b111111111111;
assign Lowerletter[792] = 12'b111111111111;
assign Lowerletter[793] = 12'b000000000000;
assign Lowerletter[794] = 12'b111111111111;
assign Lowerletter[795] = 12'b000000000000;
assign Lowerletter[796] = 12'b111111111111;
assign Lowerletter[797] = 12'b000000000000;
assign Lowerletter[798] = 12'b111111111111;
assign Lowerletter[799] = 12'b111111111111;
assign Lowerletter[800] = 12'b111111111111;
assign Lowerletter[801] = 12'b000000000000;
assign Lowerletter[802] = 12'b111111111111;
assign Lowerletter[803] = 12'b000000000000;
assign Lowerletter[804] = 12'b111111111111;
assign Lowerletter[805] = 12'b000000000000;
assign Lowerletter[806] = 12'b111111111111;
assign Lowerletter[807] = 12'b111111111111;
assign Lowerletter[808] = 12'b111111111111;
assign Lowerletter[809] = 12'b000000000000;
assign Lowerletter[810] = 12'b111111111111;
assign Lowerletter[811] = 12'b000000000000;
assign Lowerletter[812] = 12'b111111111111;
assign Lowerletter[813] = 12'b000000000000;
assign Lowerletter[814] = 12'b111111111111;
assign Lowerletter[815] = 12'b111111111111;
assign Lowerletter[816] = 12'b111111111111;
assign Lowerletter[817] = 12'b000000000000;
assign Lowerletter[818] = 12'b111111111111;
assign Lowerletter[819] = 12'b000000000000;
assign Lowerletter[820] = 12'b111111111111;
assign Lowerletter[821] = 12'b000000000000;
assign Lowerletter[822] = 12'b111111111111;
assign Lowerletter[823] = 12'b111111111111;
assign Lowerletter[824] = 12'b111111111111;
assign Lowerletter[825] = 12'b111111111111;
assign Lowerletter[826] = 12'b111111111111;
assign Lowerletter[827] = 12'b111111111111;
assign Lowerletter[828] = 12'b111111111111;
assign Lowerletter[829] = 12'b111111111111;
assign Lowerletter[830] = 12'b111111111111;
assign Lowerletter[831] = 12'b111111111111;
assign Lowerletter[832] = 12'b111111111111;
assign Lowerletter[833] = 12'b111111111111;
assign Lowerletter[834] = 12'b111111111111;
assign Lowerletter[835] = 12'b111111111111;
assign Lowerletter[836] = 12'b111111111111;
assign Lowerletter[837] = 12'b111111111111;
assign Lowerletter[838] = 12'b111111111111;
assign Lowerletter[839] = 12'b111111111111;
assign Lowerletter[840] = 12'b111111111111;
assign Lowerletter[841] = 12'b111111111111;
assign Lowerletter[842] = 12'b111111111111;
assign Lowerletter[843] = 12'b111111111111;
assign Lowerletter[844] = 12'b111111111111;
assign Lowerletter[845] = 12'b111111111111;
assign Lowerletter[846] = 12'b111111111111;
assign Lowerletter[847] = 12'b111111111111;
assign Lowerletter[848] = 12'b111111111111;
assign Lowerletter[849] = 12'b111111111111;
assign Lowerletter[850] = 12'b000000000000;
assign Lowerletter[851] = 12'b000000000000;
assign Lowerletter[852] = 12'b000000000000;
assign Lowerletter[853] = 12'b111111111111;
assign Lowerletter[854] = 12'b111111111111;
assign Lowerletter[855] = 12'b111111111111;
assign Lowerletter[856] = 12'b111111111111;
assign Lowerletter[857] = 12'b111111111111;
assign Lowerletter[858] = 12'b000000000000;
assign Lowerletter[859] = 12'b111111111111;
assign Lowerletter[860] = 12'b111111111111;
assign Lowerletter[861] = 12'b000000000000;
assign Lowerletter[862] = 12'b111111111111;
assign Lowerletter[863] = 12'b111111111111;
assign Lowerletter[864] = 12'b111111111111;
assign Lowerletter[865] = 12'b111111111111;
assign Lowerletter[866] = 12'b000000000000;
assign Lowerletter[867] = 12'b111111111111;
assign Lowerletter[868] = 12'b111111111111;
assign Lowerletter[869] = 12'b000000000000;
assign Lowerletter[870] = 12'b111111111111;
assign Lowerletter[871] = 12'b111111111111;
assign Lowerletter[872] = 12'b111111111111;
assign Lowerletter[873] = 12'b111111111111;
assign Lowerletter[874] = 12'b000000000000;
assign Lowerletter[875] = 12'b111111111111;
assign Lowerletter[876] = 12'b111111111111;
assign Lowerletter[877] = 12'b000000000000;
assign Lowerletter[878] = 12'b111111111111;
assign Lowerletter[879] = 12'b111111111111;
assign Lowerletter[880] = 12'b111111111111;
assign Lowerletter[881] = 12'b111111111111;
assign Lowerletter[882] = 12'b000000000000;
assign Lowerletter[883] = 12'b111111111111;
assign Lowerletter[884] = 12'b111111111111;
assign Lowerletter[885] = 12'b000000000000;
assign Lowerletter[886] = 12'b111111111111;
assign Lowerletter[887] = 12'b111111111111;
assign Lowerletter[888] = 12'b111111111111;
assign Lowerletter[889] = 12'b111111111111;
assign Lowerletter[890] = 12'b111111111111;
assign Lowerletter[891] = 12'b111111111111;
assign Lowerletter[892] = 12'b111111111111;
assign Lowerletter[893] = 12'b111111111111;
assign Lowerletter[894] = 12'b111111111111;
assign Lowerletter[895] = 12'b111111111111;
assign Lowerletter[896] = 12'b111111111111;
assign Lowerletter[897] = 12'b111111111111;
assign Lowerletter[898] = 12'b111111111111;
assign Lowerletter[899] = 12'b111111111111;
assign Lowerletter[900] = 12'b111111111111;
assign Lowerletter[901] = 12'b111111111111;
assign Lowerletter[902] = 12'b111111111111;
assign Lowerletter[903] = 12'b111111111111;
assign Lowerletter[904] = 12'b111111111111;
assign Lowerletter[905] = 12'b111111111111;
assign Lowerletter[906] = 12'b111111111111;
assign Lowerletter[907] = 12'b111111111111;
assign Lowerletter[908] = 12'b111111111111;
assign Lowerletter[909] = 12'b111111111111;
assign Lowerletter[910] = 12'b111111111111;
assign Lowerletter[911] = 12'b111111111111;
assign Lowerletter[912] = 12'b111111111111;
assign Lowerletter[913] = 12'b111111111111;
assign Lowerletter[914] = 12'b111111111111;
assign Lowerletter[915] = 12'b000000000000;
assign Lowerletter[916] = 12'b000000000000;
assign Lowerletter[917] = 12'b111111111111;
assign Lowerletter[918] = 12'b111111111111;
assign Lowerletter[919] = 12'b111111111111;
assign Lowerletter[920] = 12'b111111111111;
assign Lowerletter[921] = 12'b111111111111;
assign Lowerletter[922] = 12'b000000000000;
assign Lowerletter[923] = 12'b111111111111;
assign Lowerletter[924] = 12'b111111111111;
assign Lowerletter[925] = 12'b000000000000;
assign Lowerletter[926] = 12'b111111111111;
assign Lowerletter[927] = 12'b111111111111;
assign Lowerletter[928] = 12'b111111111111;
assign Lowerletter[929] = 12'b111111111111;
assign Lowerletter[930] = 12'b000000000000;
assign Lowerletter[931] = 12'b111111111111;
assign Lowerletter[932] = 12'b111111111111;
assign Lowerletter[933] = 12'b000000000000;
assign Lowerletter[934] = 12'b111111111111;
assign Lowerletter[935] = 12'b111111111111;
assign Lowerletter[936] = 12'b111111111111;
assign Lowerletter[937] = 12'b111111111111;
assign Lowerletter[938] = 12'b000000000000;
assign Lowerletter[939] = 12'b111111111111;
assign Lowerletter[940] = 12'b111111111111;
assign Lowerletter[941] = 12'b000000000000;
assign Lowerletter[942] = 12'b111111111111;
assign Lowerletter[943] = 12'b111111111111;
assign Lowerletter[944] = 12'b111111111111;
assign Lowerletter[945] = 12'b111111111111;
assign Lowerletter[946] = 12'b111111111111;
assign Lowerletter[947] = 12'b000000000000;
assign Lowerletter[948] = 12'b000000000000;
assign Lowerletter[949] = 12'b111111111111;
assign Lowerletter[950] = 12'b111111111111;
assign Lowerletter[951] = 12'b111111111111;
assign Lowerletter[952] = 12'b111111111111;
assign Lowerletter[953] = 12'b111111111111;
assign Lowerletter[954] = 12'b111111111111;
assign Lowerletter[955] = 12'b111111111111;
assign Lowerletter[956] = 12'b111111111111;
assign Lowerletter[957] = 12'b111111111111;
assign Lowerletter[958] = 12'b111111111111;
assign Lowerletter[959] = 12'b111111111111;
assign Lowerletter[960] = 12'b111111111111;
assign Lowerletter[961] = 12'b111111111111;
assign Lowerletter[962] = 12'b111111111111;
assign Lowerletter[963] = 12'b111111111111;
assign Lowerletter[964] = 12'b111111111111;
assign Lowerletter[965] = 12'b111111111111;
assign Lowerletter[966] = 12'b111111111111;
assign Lowerletter[967] = 12'b111111111111;
assign Lowerletter[968] = 12'b111111111111;
assign Lowerletter[969] = 12'b111111111111;
assign Lowerletter[970] = 12'b111111111111;
assign Lowerletter[971] = 12'b111111111111;
assign Lowerletter[972] = 12'b111111111111;
assign Lowerletter[973] = 12'b111111111111;
assign Lowerletter[974] = 12'b111111111111;
assign Lowerletter[975] = 12'b111111111111;
assign Lowerletter[976] = 12'b111111111111;
assign Lowerletter[977] = 12'b111111111111;
assign Lowerletter[978] = 12'b000000000000;
assign Lowerletter[979] = 12'b111111111111;
assign Lowerletter[980] = 12'b000000000000;
assign Lowerletter[981] = 12'b111111111111;
assign Lowerletter[982] = 12'b111111111111;
assign Lowerletter[983] = 12'b111111111111;
assign Lowerletter[984] = 12'b111111111111;
assign Lowerletter[985] = 12'b111111111111;
assign Lowerletter[986] = 12'b000000000000;
assign Lowerletter[987] = 12'b000000000000;
assign Lowerletter[988] = 12'b111111111111;
assign Lowerletter[989] = 12'b000000000000;
assign Lowerletter[990] = 12'b111111111111;
assign Lowerletter[991] = 12'b111111111111;
assign Lowerletter[992] = 12'b111111111111;
assign Lowerletter[993] = 12'b111111111111;
assign Lowerletter[994] = 12'b000000000000;
assign Lowerletter[995] = 12'b111111111111;
assign Lowerletter[996] = 12'b111111111111;
assign Lowerletter[997] = 12'b000000000000;
assign Lowerletter[998] = 12'b111111111111;
assign Lowerletter[999] = 12'b111111111111;
assign Lowerletter[1000] = 12'b111111111111;
assign Lowerletter[1001] = 12'b111111111111;
assign Lowerletter[1002] = 12'b000000000000;
assign Lowerletter[1003] = 12'b000000000000;
assign Lowerletter[1004] = 12'b000000000000;
assign Lowerletter[1005] = 12'b111111111111;
assign Lowerletter[1006] = 12'b111111111111;
assign Lowerletter[1007] = 12'b111111111111;
assign Lowerletter[1008] = 12'b111111111111;
assign Lowerletter[1009] = 12'b111111111111;
assign Lowerletter[1010] = 12'b000000000000;
assign Lowerletter[1011] = 12'b111111111111;
assign Lowerletter[1012] = 12'b111111111111;
assign Lowerletter[1013] = 12'b111111111111;
assign Lowerletter[1014] = 12'b111111111111;
assign Lowerletter[1015] = 12'b111111111111;
assign Lowerletter[1016] = 12'b111111111111;
assign Lowerletter[1017] = 12'b111111111111;
assign Lowerletter[1018] = 12'b000000000000;
assign Lowerletter[1019] = 12'b111111111111;
assign Lowerletter[1020] = 12'b111111111111;
assign Lowerletter[1021] = 12'b111111111111;
assign Lowerletter[1022] = 12'b111111111111;
assign Lowerletter[1023] = 12'b111111111111;
assign Lowerletter[1024] = 12'b111111111111;
assign Lowerletter[1025] = 12'b111111111111;
assign Lowerletter[1026] = 12'b111111111111;
assign Lowerletter[1027] = 12'b111111111111;
assign Lowerletter[1028] = 12'b111111111111;
assign Lowerletter[1029] = 12'b111111111111;
assign Lowerletter[1030] = 12'b111111111111;
assign Lowerletter[1031] = 12'b111111111111;
assign Lowerletter[1032] = 12'b111111111111;
assign Lowerletter[1033] = 12'b111111111111;
assign Lowerletter[1034] = 12'b111111111111;
assign Lowerletter[1035] = 12'b111111111111;
assign Lowerletter[1036] = 12'b111111111111;
assign Lowerletter[1037] = 12'b111111111111;
assign Lowerletter[1038] = 12'b111111111111;
assign Lowerletter[1039] = 12'b111111111111;
assign Lowerletter[1040] = 12'b111111111111;
assign Lowerletter[1041] = 12'b111111111111;
assign Lowerletter[1042] = 12'b111111111111;
assign Lowerletter[1043] = 12'b000000000000;
assign Lowerletter[1044] = 12'b111111111111;
assign Lowerletter[1045] = 12'b000000000000;
assign Lowerletter[1046] = 12'b111111111111;
assign Lowerletter[1047] = 12'b111111111111;
assign Lowerletter[1048] = 12'b111111111111;
assign Lowerletter[1049] = 12'b111111111111;
assign Lowerletter[1050] = 12'b000000000000;
assign Lowerletter[1051] = 12'b111111111111;
assign Lowerletter[1052] = 12'b000000000000;
assign Lowerletter[1053] = 12'b000000000000;
assign Lowerletter[1054] = 12'b111111111111;
assign Lowerletter[1055] = 12'b111111111111;
assign Lowerletter[1056] = 12'b111111111111;
assign Lowerletter[1057] = 12'b111111111111;
assign Lowerletter[1058] = 12'b000000000000;
assign Lowerletter[1059] = 12'b111111111111;
assign Lowerletter[1060] = 12'b111111111111;
assign Lowerletter[1061] = 12'b000000000000;
assign Lowerletter[1062] = 12'b111111111111;
assign Lowerletter[1063] = 12'b111111111111;
assign Lowerletter[1064] = 12'b111111111111;
assign Lowerletter[1065] = 12'b111111111111;
assign Lowerletter[1066] = 12'b111111111111;
assign Lowerletter[1067] = 12'b000000000000;
assign Lowerletter[1068] = 12'b000000000000;
assign Lowerletter[1069] = 12'b000000000000;
assign Lowerletter[1070] = 12'b111111111111;
assign Lowerletter[1071] = 12'b111111111111;
assign Lowerletter[1072] = 12'b111111111111;
assign Lowerletter[1073] = 12'b111111111111;
assign Lowerletter[1074] = 12'b111111111111;
assign Lowerletter[1075] = 12'b111111111111;
assign Lowerletter[1076] = 12'b111111111111;
assign Lowerletter[1077] = 12'b000000000000;
assign Lowerletter[1078] = 12'b111111111111;
assign Lowerletter[1079] = 12'b111111111111;
assign Lowerletter[1080] = 12'b111111111111;
assign Lowerletter[1081] = 12'b111111111111;
assign Lowerletter[1082] = 12'b111111111111;
assign Lowerletter[1083] = 12'b111111111111;
assign Lowerletter[1084] = 12'b111111111111;
assign Lowerletter[1085] = 12'b000000000000;
assign Lowerletter[1086] = 12'b111111111111;
assign Lowerletter[1087] = 12'b111111111111;
assign Lowerletter[1088] = 12'b111111111111;
assign Lowerletter[1089] = 12'b111111111111;
assign Lowerletter[1090] = 12'b111111111111;
assign Lowerletter[1091] = 12'b111111111111;
assign Lowerletter[1092] = 12'b111111111111;
assign Lowerletter[1093] = 12'b111111111111;
assign Lowerletter[1094] = 12'b111111111111;
assign Lowerletter[1095] = 12'b111111111111;
assign Lowerletter[1096] = 12'b111111111111;
assign Lowerletter[1097] = 12'b111111111111;
assign Lowerletter[1098] = 12'b111111111111;
assign Lowerletter[1099] = 12'b111111111111;
assign Lowerletter[1100] = 12'b111111111111;
assign Lowerletter[1101] = 12'b111111111111;
assign Lowerletter[1102] = 12'b111111111111;
assign Lowerletter[1103] = 12'b111111111111;
assign Lowerletter[1104] = 12'b111111111111;
assign Lowerletter[1105] = 12'b111111111111;
assign Lowerletter[1106] = 12'b000000000000;
assign Lowerletter[1107] = 12'b111111111111;
assign Lowerletter[1108] = 12'b000000000000;
assign Lowerletter[1109] = 12'b000000000000;
assign Lowerletter[1110] = 12'b111111111111;
assign Lowerletter[1111] = 12'b111111111111;
assign Lowerletter[1112] = 12'b111111111111;
assign Lowerletter[1113] = 12'b111111111111;
assign Lowerletter[1114] = 12'b000000000000;
assign Lowerletter[1115] = 12'b000000000000;
assign Lowerletter[1116] = 12'b111111111111;
assign Lowerletter[1117] = 12'b111111111111;
assign Lowerletter[1118] = 12'b111111111111;
assign Lowerletter[1119] = 12'b111111111111;
assign Lowerletter[1120] = 12'b111111111111;
assign Lowerletter[1121] = 12'b111111111111;
assign Lowerletter[1122] = 12'b000000000000;
assign Lowerletter[1123] = 12'b111111111111;
assign Lowerletter[1124] = 12'b111111111111;
assign Lowerletter[1125] = 12'b111111111111;
assign Lowerletter[1126] = 12'b111111111111;
assign Lowerletter[1127] = 12'b111111111111;
assign Lowerletter[1128] = 12'b111111111111;
assign Lowerletter[1129] = 12'b111111111111;
assign Lowerletter[1130] = 12'b000000000000;
assign Lowerletter[1131] = 12'b111111111111;
assign Lowerletter[1132] = 12'b111111111111;
assign Lowerletter[1133] = 12'b111111111111;
assign Lowerletter[1134] = 12'b111111111111;
assign Lowerletter[1135] = 12'b111111111111;
assign Lowerletter[1136] = 12'b111111111111;
assign Lowerletter[1137] = 12'b111111111111;
assign Lowerletter[1138] = 12'b000000000000;
assign Lowerletter[1139] = 12'b111111111111;
assign Lowerletter[1140] = 12'b111111111111;
assign Lowerletter[1141] = 12'b111111111111;
assign Lowerletter[1142] = 12'b111111111111;
assign Lowerletter[1143] = 12'b111111111111;
assign Lowerletter[1144] = 12'b111111111111;
assign Lowerletter[1145] = 12'b111111111111;
assign Lowerletter[1146] = 12'b111111111111;
assign Lowerletter[1147] = 12'b111111111111;
assign Lowerletter[1148] = 12'b111111111111;
assign Lowerletter[1149] = 12'b111111111111;
assign Lowerletter[1150] = 12'b111111111111;
assign Lowerletter[1151] = 12'b111111111111;
assign Lowerletter[1152] = 12'b111111111111;
assign Lowerletter[1153] = 12'b111111111111;
assign Lowerletter[1154] = 12'b111111111111;
assign Lowerletter[1155] = 12'b111111111111;
assign Lowerletter[1156] = 12'b111111111111;
assign Lowerletter[1157] = 12'b111111111111;
assign Lowerletter[1158] = 12'b111111111111;
assign Lowerletter[1159] = 12'b111111111111;
assign Lowerletter[1160] = 12'b111111111111;
assign Lowerletter[1161] = 12'b111111111111;
assign Lowerletter[1162] = 12'b111111111111;
assign Lowerletter[1163] = 12'b111111111111;
assign Lowerletter[1164] = 12'b111111111111;
assign Lowerletter[1165] = 12'b111111111111;
assign Lowerletter[1166] = 12'b111111111111;
assign Lowerletter[1167] = 12'b111111111111;
assign Lowerletter[1168] = 12'b111111111111;
assign Lowerletter[1169] = 12'b111111111111;
assign Lowerletter[1170] = 12'b111111111111;
assign Lowerletter[1171] = 12'b000000000000;
assign Lowerletter[1172] = 12'b000000000000;
assign Lowerletter[1173] = 12'b000000000000;
assign Lowerletter[1174] = 12'b111111111111;
assign Lowerletter[1175] = 12'b111111111111;
assign Lowerletter[1176] = 12'b111111111111;
assign Lowerletter[1177] = 12'b111111111111;
assign Lowerletter[1178] = 12'b000000000000;
assign Lowerletter[1179] = 12'b111111111111;
assign Lowerletter[1180] = 12'b111111111111;
assign Lowerletter[1181] = 12'b111111111111;
assign Lowerletter[1182] = 12'b111111111111;
assign Lowerletter[1183] = 12'b111111111111;
assign Lowerletter[1184] = 12'b111111111111;
assign Lowerletter[1185] = 12'b111111111111;
assign Lowerletter[1186] = 12'b111111111111;
assign Lowerletter[1187] = 12'b000000000000;
assign Lowerletter[1188] = 12'b000000000000;
assign Lowerletter[1189] = 12'b111111111111;
assign Lowerletter[1190] = 12'b111111111111;
assign Lowerletter[1191] = 12'b111111111111;
assign Lowerletter[1192] = 12'b111111111111;
assign Lowerletter[1193] = 12'b111111111111;
assign Lowerletter[1194] = 12'b111111111111;
assign Lowerletter[1195] = 12'b111111111111;
assign Lowerletter[1196] = 12'b111111111111;
assign Lowerletter[1197] = 12'b000000000000;
assign Lowerletter[1198] = 12'b111111111111;
assign Lowerletter[1199] = 12'b111111111111;
assign Lowerletter[1200] = 12'b111111111111;
assign Lowerletter[1201] = 12'b111111111111;
assign Lowerletter[1202] = 12'b000000000000;
assign Lowerletter[1203] = 12'b000000000000;
assign Lowerletter[1204] = 12'b000000000000;
assign Lowerletter[1205] = 12'b111111111111;
assign Lowerletter[1206] = 12'b111111111111;
assign Lowerletter[1207] = 12'b111111111111;
assign Lowerletter[1208] = 12'b111111111111;
assign Lowerletter[1209] = 12'b111111111111;
assign Lowerletter[1210] = 12'b111111111111;
assign Lowerletter[1211] = 12'b111111111111;
assign Lowerletter[1212] = 12'b111111111111;
assign Lowerletter[1213] = 12'b111111111111;
assign Lowerletter[1214] = 12'b111111111111;
assign Lowerletter[1215] = 12'b111111111111;
assign Lowerletter[1216] = 12'b111111111111;
assign Lowerletter[1217] = 12'b111111111111;
assign Lowerletter[1218] = 12'b111111111111;
assign Lowerletter[1219] = 12'b111111111111;
assign Lowerletter[1220] = 12'b111111111111;
assign Lowerletter[1221] = 12'b111111111111;
assign Lowerletter[1222] = 12'b111111111111;
assign Lowerletter[1223] = 12'b111111111111;
assign Lowerletter[1224] = 12'b111111111111;
assign Lowerletter[1225] = 12'b111111111111;
assign Lowerletter[1226] = 12'b111111111111;
assign Lowerletter[1227] = 12'b000000000000;
assign Lowerletter[1228] = 12'b111111111111;
assign Lowerletter[1229] = 12'b111111111111;
assign Lowerletter[1230] = 12'b111111111111;
assign Lowerletter[1231] = 12'b111111111111;
assign Lowerletter[1232] = 12'b111111111111;
assign Lowerletter[1233] = 12'b111111111111;
assign Lowerletter[1234] = 12'b000000000000;
assign Lowerletter[1235] = 12'b000000000000;
assign Lowerletter[1236] = 12'b000000000000;
assign Lowerletter[1237] = 12'b111111111111;
assign Lowerletter[1238] = 12'b111111111111;
assign Lowerletter[1239] = 12'b111111111111;
assign Lowerletter[1240] = 12'b111111111111;
assign Lowerletter[1241] = 12'b111111111111;
assign Lowerletter[1242] = 12'b111111111111;
assign Lowerletter[1243] = 12'b000000000000;
assign Lowerletter[1244] = 12'b111111111111;
assign Lowerletter[1245] = 12'b111111111111;
assign Lowerletter[1246] = 12'b111111111111;
assign Lowerletter[1247] = 12'b111111111111;
assign Lowerletter[1248] = 12'b111111111111;
assign Lowerletter[1249] = 12'b111111111111;
assign Lowerletter[1250] = 12'b111111111111;
assign Lowerletter[1251] = 12'b000000000000;
assign Lowerletter[1252] = 12'b111111111111;
assign Lowerletter[1253] = 12'b111111111111;
assign Lowerletter[1254] = 12'b111111111111;
assign Lowerletter[1255] = 12'b111111111111;
assign Lowerletter[1256] = 12'b111111111111;
assign Lowerletter[1257] = 12'b111111111111;
assign Lowerletter[1258] = 12'b111111111111;
assign Lowerletter[1259] = 12'b000000000000;
assign Lowerletter[1260] = 12'b111111111111;
assign Lowerletter[1261] = 12'b111111111111;
assign Lowerletter[1262] = 12'b111111111111;
assign Lowerletter[1263] = 12'b111111111111;
assign Lowerletter[1264] = 12'b111111111111;
assign Lowerletter[1265] = 12'b111111111111;
assign Lowerletter[1266] = 12'b111111111111;
assign Lowerletter[1267] = 12'b111111111111;
assign Lowerletter[1268] = 12'b000000000000;
assign Lowerletter[1269] = 12'b111111111111;
assign Lowerletter[1270] = 12'b111111111111;
assign Lowerletter[1271] = 12'b111111111111;
assign Lowerletter[1272] = 12'b111111111111;
assign Lowerletter[1273] = 12'b111111111111;
assign Lowerletter[1274] = 12'b111111111111;
assign Lowerletter[1275] = 12'b111111111111;
assign Lowerletter[1276] = 12'b111111111111;
assign Lowerletter[1277] = 12'b111111111111;
assign Lowerletter[1278] = 12'b111111111111;
assign Lowerletter[1279] = 12'b111111111111;
assign Lowerletter[1280] = 12'b111111111111;
assign Lowerletter[1281] = 12'b111111111111;
assign Lowerletter[1282] = 12'b111111111111;
assign Lowerletter[1283] = 12'b111111111111;
assign Lowerletter[1284] = 12'b111111111111;
assign Lowerletter[1285] = 12'b111111111111;
assign Lowerletter[1286] = 12'b111111111111;
assign Lowerletter[1287] = 12'b111111111111;
assign Lowerletter[1288] = 12'b111111111111;
assign Lowerletter[1289] = 12'b111111111111;
assign Lowerletter[1290] = 12'b111111111111;
assign Lowerletter[1291] = 12'b111111111111;
assign Lowerletter[1292] = 12'b111111111111;
assign Lowerletter[1293] = 12'b111111111111;
assign Lowerletter[1294] = 12'b111111111111;
assign Lowerletter[1295] = 12'b111111111111;
assign Lowerletter[1296] = 12'b111111111111;
assign Lowerletter[1297] = 12'b111111111111;
assign Lowerletter[1298] = 12'b000000000000;
assign Lowerletter[1299] = 12'b111111111111;
assign Lowerletter[1300] = 12'b111111111111;
assign Lowerletter[1301] = 12'b000000000000;
assign Lowerletter[1302] = 12'b111111111111;
assign Lowerletter[1303] = 12'b111111111111;
assign Lowerletter[1304] = 12'b111111111111;
assign Lowerletter[1305] = 12'b111111111111;
assign Lowerletter[1306] = 12'b000000000000;
assign Lowerletter[1307] = 12'b111111111111;
assign Lowerletter[1308] = 12'b111111111111;
assign Lowerletter[1309] = 12'b000000000000;
assign Lowerletter[1310] = 12'b111111111111;
assign Lowerletter[1311] = 12'b111111111111;
assign Lowerletter[1312] = 12'b111111111111;
assign Lowerletter[1313] = 12'b111111111111;
assign Lowerletter[1314] = 12'b000000000000;
assign Lowerletter[1315] = 12'b111111111111;
assign Lowerletter[1316] = 12'b111111111111;
assign Lowerletter[1317] = 12'b000000000000;
assign Lowerletter[1318] = 12'b111111111111;
assign Lowerletter[1319] = 12'b111111111111;
assign Lowerletter[1320] = 12'b111111111111;
assign Lowerletter[1321] = 12'b111111111111;
assign Lowerletter[1322] = 12'b000000000000;
assign Lowerletter[1323] = 12'b111111111111;
assign Lowerletter[1324] = 12'b111111111111;
assign Lowerletter[1325] = 12'b000000000000;
assign Lowerletter[1326] = 12'b111111111111;
assign Lowerletter[1327] = 12'b111111111111;
assign Lowerletter[1328] = 12'b111111111111;
assign Lowerletter[1329] = 12'b111111111111;
assign Lowerletter[1330] = 12'b111111111111;
assign Lowerletter[1331] = 12'b000000000000;
assign Lowerletter[1332] = 12'b000000000000;
assign Lowerletter[1333] = 12'b111111111111;
assign Lowerletter[1334] = 12'b111111111111;
assign Lowerletter[1335] = 12'b111111111111;
assign Lowerletter[1336] = 12'b111111111111;
assign Lowerletter[1337] = 12'b111111111111;
assign Lowerletter[1338] = 12'b111111111111;
assign Lowerletter[1339] = 12'b111111111111;
assign Lowerletter[1340] = 12'b111111111111;
assign Lowerletter[1341] = 12'b111111111111;
assign Lowerletter[1342] = 12'b111111111111;
assign Lowerletter[1343] = 12'b111111111111;
assign Lowerletter[1344] = 12'b111111111111;
assign Lowerletter[1345] = 12'b111111111111;
assign Lowerletter[1346] = 12'b111111111111;
assign Lowerletter[1347] = 12'b111111111111;
assign Lowerletter[1348] = 12'b111111111111;
assign Lowerletter[1349] = 12'b111111111111;
assign Lowerletter[1350] = 12'b111111111111;
assign Lowerletter[1351] = 12'b111111111111;
assign Lowerletter[1352] = 12'b111111111111;
assign Lowerletter[1353] = 12'b111111111111;
assign Lowerletter[1354] = 12'b111111111111;
assign Lowerletter[1355] = 12'b111111111111;
assign Lowerletter[1356] = 12'b111111111111;
assign Lowerletter[1357] = 12'b111111111111;
assign Lowerletter[1358] = 12'b111111111111;
assign Lowerletter[1359] = 12'b111111111111;
assign Lowerletter[1360] = 12'b111111111111;
assign Lowerletter[1361] = 12'b000000000000;
assign Lowerletter[1362] = 12'b111111111111;
assign Lowerletter[1363] = 12'b111111111111;
assign Lowerletter[1364] = 12'b111111111111;
assign Lowerletter[1365] = 12'b000000000000;
assign Lowerletter[1366] = 12'b111111111111;
assign Lowerletter[1367] = 12'b111111111111;
assign Lowerletter[1368] = 12'b111111111111;
assign Lowerletter[1369] = 12'b000000000000;
assign Lowerletter[1370] = 12'b111111111111;
assign Lowerletter[1371] = 12'b111111111111;
assign Lowerletter[1372] = 12'b111111111111;
assign Lowerletter[1373] = 12'b000000000000;
assign Lowerletter[1374] = 12'b111111111111;
assign Lowerletter[1375] = 12'b111111111111;
assign Lowerletter[1376] = 12'b111111111111;
assign Lowerletter[1377] = 12'b000000000000;
assign Lowerletter[1378] = 12'b111111111111;
assign Lowerletter[1379] = 12'b111111111111;
assign Lowerletter[1380] = 12'b111111111111;
assign Lowerletter[1381] = 12'b000000000000;
assign Lowerletter[1382] = 12'b111111111111;
assign Lowerletter[1383] = 12'b111111111111;
assign Lowerletter[1384] = 12'b111111111111;
assign Lowerletter[1385] = 12'b111111111111;
assign Lowerletter[1386] = 12'b000000000000;
assign Lowerletter[1387] = 12'b111111111111;
assign Lowerletter[1388] = 12'b000000000000;
assign Lowerletter[1389] = 12'b111111111111;
assign Lowerletter[1390] = 12'b111111111111;
assign Lowerletter[1391] = 12'b111111111111;
assign Lowerletter[1392] = 12'b111111111111;
assign Lowerletter[1393] = 12'b111111111111;
assign Lowerletter[1394] = 12'b111111111111;
assign Lowerletter[1395] = 12'b000000000000;
assign Lowerletter[1396] = 12'b111111111111;
assign Lowerletter[1397] = 12'b111111111111;
assign Lowerletter[1398] = 12'b111111111111;
assign Lowerletter[1399] = 12'b111111111111;
assign Lowerletter[1400] = 12'b111111111111;
assign Lowerletter[1401] = 12'b111111111111;
assign Lowerletter[1402] = 12'b111111111111;
assign Lowerletter[1403] = 12'b111111111111;
assign Lowerletter[1404] = 12'b111111111111;
assign Lowerletter[1405] = 12'b111111111111;
assign Lowerletter[1406] = 12'b111111111111;
assign Lowerletter[1407] = 12'b111111111111;
assign Lowerletter[1408] = 12'b111111111111;
assign Lowerletter[1409] = 12'b111111111111;
assign Lowerletter[1410] = 12'b111111111111;
assign Lowerletter[1411] = 12'b111111111111;
assign Lowerletter[1412] = 12'b111111111111;
assign Lowerletter[1413] = 12'b111111111111;
assign Lowerletter[1414] = 12'b111111111111;
assign Lowerletter[1415] = 12'b111111111111;
assign Lowerletter[1416] = 12'b111111111111;
assign Lowerletter[1417] = 12'b111111111111;
assign Lowerletter[1418] = 12'b111111111111;
assign Lowerletter[1419] = 12'b111111111111;
assign Lowerletter[1420] = 12'b111111111111;
assign Lowerletter[1421] = 12'b111111111111;
assign Lowerletter[1422] = 12'b111111111111;
assign Lowerletter[1423] = 12'b111111111111;
assign Lowerletter[1424] = 12'b111111111111;
assign Lowerletter[1425] = 12'b111111111111;
assign Lowerletter[1426] = 12'b111111111111;
assign Lowerletter[1427] = 12'b111111111111;
assign Lowerletter[1428] = 12'b111111111111;
assign Lowerletter[1429] = 12'b111111111111;
assign Lowerletter[1430] = 12'b111111111111;
assign Lowerletter[1431] = 12'b111111111111;
assign Lowerletter[1432] = 12'b111111111111;
assign Lowerletter[1433] = 12'b000000000000;
assign Lowerletter[1434] = 12'b111111111111;
assign Lowerletter[1435] = 12'b111111111111;
assign Lowerletter[1436] = 12'b111111111111;
assign Lowerletter[1437] = 12'b000000000000;
assign Lowerletter[1438] = 12'b111111111111;
assign Lowerletter[1439] = 12'b111111111111;
assign Lowerletter[1440] = 12'b111111111111;
assign Lowerletter[1441] = 12'b000000000000;
assign Lowerletter[1442] = 12'b111111111111;
assign Lowerletter[1443] = 12'b111111111111;
assign Lowerletter[1444] = 12'b111111111111;
assign Lowerletter[1445] = 12'b000000000000;
assign Lowerletter[1446] = 12'b111111111111;
assign Lowerletter[1447] = 12'b111111111111;
assign Lowerletter[1448] = 12'b111111111111;
assign Lowerletter[1449] = 12'b000000000000;
assign Lowerletter[1450] = 12'b111111111111;
assign Lowerletter[1451] = 12'b000000000000;
assign Lowerletter[1452] = 12'b111111111111;
assign Lowerletter[1453] = 12'b000000000000;
assign Lowerletter[1454] = 12'b111111111111;
assign Lowerletter[1455] = 12'b111111111111;
assign Lowerletter[1456] = 12'b111111111111;
assign Lowerletter[1457] = 12'b111111111111;
assign Lowerletter[1458] = 12'b000000000000;
assign Lowerletter[1459] = 12'b000000000000;
assign Lowerletter[1460] = 12'b000000000000;
assign Lowerletter[1461] = 12'b000000000000;
assign Lowerletter[1462] = 12'b111111111111;
assign Lowerletter[1463] = 12'b111111111111;
assign Lowerletter[1464] = 12'b111111111111;
assign Lowerletter[1465] = 12'b111111111111;
assign Lowerletter[1466] = 12'b111111111111;
assign Lowerletter[1467] = 12'b111111111111;
assign Lowerletter[1468] = 12'b111111111111;
assign Lowerletter[1469] = 12'b111111111111;
assign Lowerletter[1470] = 12'b111111111111;
assign Lowerletter[1471] = 12'b111111111111;
assign Lowerletter[1472] = 12'b111111111111;
assign Lowerletter[1473] = 12'b111111111111;
assign Lowerletter[1474] = 12'b111111111111;
assign Lowerletter[1475] = 12'b111111111111;
assign Lowerletter[1476] = 12'b111111111111;
assign Lowerletter[1477] = 12'b111111111111;
assign Lowerletter[1478] = 12'b111111111111;
assign Lowerletter[1479] = 12'b111111111111;
assign Lowerletter[1480] = 12'b111111111111;
assign Lowerletter[1481] = 12'b111111111111;
assign Lowerletter[1482] = 12'b111111111111;
assign Lowerletter[1483] = 12'b111111111111;
assign Lowerletter[1484] = 12'b111111111111;
assign Lowerletter[1485] = 12'b111111111111;
assign Lowerletter[1486] = 12'b111111111111;
assign Lowerletter[1487] = 12'b111111111111;
assign Lowerletter[1488] = 12'b111111111111;
assign Lowerletter[1489] = 12'b000000000000;
assign Lowerletter[1490] = 12'b111111111111;
assign Lowerletter[1491] = 12'b111111111111;
assign Lowerletter[1492] = 12'b111111111111;
assign Lowerletter[1493] = 12'b000000000000;
assign Lowerletter[1494] = 12'b111111111111;
assign Lowerletter[1495] = 12'b111111111111;
assign Lowerletter[1496] = 12'b111111111111;
assign Lowerletter[1497] = 12'b111111111111;
assign Lowerletter[1498] = 12'b000000000000;
assign Lowerletter[1499] = 12'b111111111111;
assign Lowerletter[1500] = 12'b000000000000;
assign Lowerletter[1501] = 12'b111111111111;
assign Lowerletter[1502] = 12'b111111111111;
assign Lowerletter[1503] = 12'b111111111111;
assign Lowerletter[1504] = 12'b111111111111;
assign Lowerletter[1505] = 12'b111111111111;
assign Lowerletter[1506] = 12'b111111111111;
assign Lowerletter[1507] = 12'b000000000000;
assign Lowerletter[1508] = 12'b111111111111;
assign Lowerletter[1509] = 12'b111111111111;
assign Lowerletter[1510] = 12'b111111111111;
assign Lowerletter[1511] = 12'b111111111111;
assign Lowerletter[1512] = 12'b111111111111;
assign Lowerletter[1513] = 12'b111111111111;
assign Lowerletter[1514] = 12'b000000000000;
assign Lowerletter[1515] = 12'b111111111111;
assign Lowerletter[1516] = 12'b000000000000;
assign Lowerletter[1517] = 12'b111111111111;
assign Lowerletter[1518] = 12'b111111111111;
assign Lowerletter[1519] = 12'b111111111111;
assign Lowerletter[1520] = 12'b111111111111;
assign Lowerletter[1521] = 12'b000000000000;
assign Lowerletter[1522] = 12'b111111111111;
assign Lowerletter[1523] = 12'b111111111111;
assign Lowerletter[1524] = 12'b111111111111;
assign Lowerletter[1525] = 12'b000000000000;
assign Lowerletter[1526] = 12'b111111111111;
assign Lowerletter[1527] = 12'b111111111111;
assign Lowerletter[1528] = 12'b111111111111;
assign Lowerletter[1529] = 12'b111111111111;
assign Lowerletter[1530] = 12'b111111111111;
assign Lowerletter[1531] = 12'b111111111111;
assign Lowerletter[1532] = 12'b111111111111;
assign Lowerletter[1533] = 12'b111111111111;
assign Lowerletter[1534] = 12'b111111111111;
assign Lowerletter[1535] = 12'b111111111111;
assign Lowerletter[1536] = 12'b111111111111;
assign Lowerletter[1537] = 12'b111111111111;
assign Lowerletter[1538] = 12'b111111111111;
assign Lowerletter[1539] = 12'b111111111111;
assign Lowerletter[1540] = 12'b111111111111;
assign Lowerletter[1541] = 12'b111111111111;
assign Lowerletter[1542] = 12'b111111111111;
assign Lowerletter[1543] = 12'b111111111111;
assign Lowerletter[1544] = 12'b111111111111;
assign Lowerletter[1545] = 12'b111111111111;
assign Lowerletter[1546] = 12'b111111111111;
assign Lowerletter[1547] = 12'b111111111111;
assign Lowerletter[1548] = 12'b111111111111;
assign Lowerletter[1549] = 12'b111111111111;
assign Lowerletter[1550] = 12'b111111111111;
assign Lowerletter[1551] = 12'b111111111111;
assign Lowerletter[1552] = 12'b111111111111;
assign Lowerletter[1553] = 12'b111111111111;
assign Lowerletter[1554] = 12'b000000000000;
assign Lowerletter[1555] = 12'b111111111111;
assign Lowerletter[1556] = 12'b111111111111;
assign Lowerletter[1557] = 12'b000000000000;
assign Lowerletter[1558] = 12'b111111111111;
assign Lowerletter[1559] = 12'b111111111111;
assign Lowerletter[1560] = 12'b111111111111;
assign Lowerletter[1561] = 12'b111111111111;
assign Lowerletter[1562] = 12'b000000000000;
assign Lowerletter[1563] = 12'b111111111111;
assign Lowerletter[1564] = 12'b111111111111;
assign Lowerletter[1565] = 12'b000000000000;
assign Lowerletter[1566] = 12'b111111111111;
assign Lowerletter[1567] = 12'b111111111111;
assign Lowerletter[1568] = 12'b111111111111;
assign Lowerletter[1569] = 12'b111111111111;
assign Lowerletter[1570] = 12'b000000000000;
assign Lowerletter[1571] = 12'b111111111111;
assign Lowerletter[1572] = 12'b111111111111;
assign Lowerletter[1573] = 12'b000000000000;
assign Lowerletter[1574] = 12'b111111111111;
assign Lowerletter[1575] = 12'b111111111111;
assign Lowerletter[1576] = 12'b111111111111;
assign Lowerletter[1577] = 12'b111111111111;
assign Lowerletter[1578] = 12'b111111111111;
assign Lowerletter[1579] = 12'b000000000000;
assign Lowerletter[1580] = 12'b000000000000;
assign Lowerletter[1581] = 12'b000000000000;
assign Lowerletter[1582] = 12'b111111111111;
assign Lowerletter[1583] = 12'b111111111111;
assign Lowerletter[1584] = 12'b111111111111;
assign Lowerletter[1585] = 12'b111111111111;
assign Lowerletter[1586] = 12'b111111111111;
assign Lowerletter[1587] = 12'b111111111111;
assign Lowerletter[1588] = 12'b111111111111;
assign Lowerletter[1589] = 12'b000000000000;
assign Lowerletter[1590] = 12'b111111111111;
assign Lowerletter[1591] = 12'b111111111111;
assign Lowerletter[1592] = 12'b111111111111;
assign Lowerletter[1593] = 12'b111111111111;
assign Lowerletter[1594] = 12'b000000000000;
assign Lowerletter[1595] = 12'b000000000000;
assign Lowerletter[1596] = 12'b000000000000;
assign Lowerletter[1597] = 12'b111111111111;
assign Lowerletter[1598] = 12'b111111111111;
assign Lowerletter[1599] = 12'b111111111111;
assign Lowerletter[1600] = 12'b111111111111;
assign Lowerletter[1601] = 12'b111111111111;
assign Lowerletter[1602] = 12'b111111111111;
assign Lowerletter[1603] = 12'b111111111111;
assign Lowerletter[1604] = 12'b111111111111;
assign Lowerletter[1605] = 12'b111111111111;
assign Lowerletter[1606] = 12'b111111111111;
assign Lowerletter[1607] = 12'b111111111111;
assign Lowerletter[1608] = 12'b111111111111;
assign Lowerletter[1609] = 12'b111111111111;
assign Lowerletter[1610] = 12'b111111111111;
assign Lowerletter[1611] = 12'b111111111111;
assign Lowerletter[1612] = 12'b111111111111;
assign Lowerletter[1613] = 12'b111111111111;
assign Lowerletter[1614] = 12'b111111111111;
assign Lowerletter[1615] = 12'b111111111111;
assign Lowerletter[1616] = 12'b111111111111;
assign Lowerletter[1617] = 12'b000000000000;
assign Lowerletter[1618] = 12'b000000000000;
assign Lowerletter[1619] = 12'b000000000000;
assign Lowerletter[1620] = 12'b000000000000;
assign Lowerletter[1621] = 12'b000000000000;
assign Lowerletter[1622] = 12'b111111111111;
assign Lowerletter[1623] = 12'b111111111111;
assign Lowerletter[1624] = 12'b111111111111;
assign Lowerletter[1625] = 12'b111111111111;
assign Lowerletter[1626] = 12'b111111111111;
assign Lowerletter[1627] = 12'b111111111111;
assign Lowerletter[1628] = 12'b000000000000;
assign Lowerletter[1629] = 12'b111111111111;
assign Lowerletter[1630] = 12'b111111111111;
assign Lowerletter[1631] = 12'b111111111111;
assign Lowerletter[1632] = 12'b111111111111;
assign Lowerletter[1633] = 12'b111111111111;
assign Lowerletter[1634] = 12'b111111111111;
assign Lowerletter[1635] = 12'b000000000000;
assign Lowerletter[1636] = 12'b111111111111;
assign Lowerletter[1637] = 12'b111111111111;
assign Lowerletter[1638] = 12'b111111111111;
assign Lowerletter[1639] = 12'b111111111111;
assign Lowerletter[1640] = 12'b111111111111;
assign Lowerletter[1641] = 12'b111111111111;
assign Lowerletter[1642] = 12'b000000000000;
assign Lowerletter[1643] = 12'b111111111111;
assign Lowerletter[1644] = 12'b111111111111;
assign Lowerletter[1645] = 12'b111111111111;
assign Lowerletter[1646] = 12'b111111111111;
assign Lowerletter[1647] = 12'b111111111111;
assign Lowerletter[1648] = 12'b111111111111;
assign Lowerletter[1649] = 12'b000000000000;
assign Lowerletter[1650] = 12'b000000000000;
assign Lowerletter[1651] = 12'b000000000000;
assign Lowerletter[1652] = 12'b000000000000;
assign Lowerletter[1653] = 12'b000000000000;
assign Lowerletter[1654] = 12'b111111111111;
assign Lowerletter[1655] = 12'b111111111111;
assign Lowerletter[1656] = 12'b111111111111;
assign Lowerletter[1657] = 12'b111111111111;
assign Lowerletter[1658] = 12'b111111111111;
assign Lowerletter[1659] = 12'b111111111111;
assign Lowerletter[1660] = 12'b111111111111;
assign Lowerletter[1661] = 12'b111111111111;
assign Lowerletter[1662] = 12'b111111111111;
assign Lowerletter[1663] = 12'b111111111111;
assign Upperletter[0] = 12'b111111111111;
assign Upperletter[1] = 12'b111111111111;
assign Upperletter[2] = 12'b000000000000;
assign Upperletter[3] = 12'b000000000000;
assign Upperletter[4] = 12'b000000000000;
assign Upperletter[5] = 12'b111111111111;
assign Upperletter[6] = 12'b111111111111;
assign Upperletter[7] = 12'b111111111111;
assign Upperletter[8] = 12'b111111111111;
assign Upperletter[9] = 12'b000000000000;
assign Upperletter[10] = 12'b111111111111;
assign Upperletter[11] = 12'b111111111111;
assign Upperletter[12] = 12'b111111111111;
assign Upperletter[13] = 12'b000000000000;
assign Upperletter[14] = 12'b111111111111;
assign Upperletter[15] = 12'b111111111111;
assign Upperletter[16] = 12'b111111111111;
assign Upperletter[17] = 12'b000000000000;
assign Upperletter[18] = 12'b111111111111;
assign Upperletter[19] = 12'b111111111111;
assign Upperletter[20] = 12'b111111111111;
assign Upperletter[21] = 12'b000000000000;
assign Upperletter[22] = 12'b111111111111;
assign Upperletter[23] = 12'b111111111111;
assign Upperletter[24] = 12'b111111111111;
assign Upperletter[25] = 12'b000000000000;
assign Upperletter[26] = 12'b000000000000;
assign Upperletter[27] = 12'b000000000000;
assign Upperletter[28] = 12'b000000000000;
assign Upperletter[29] = 12'b000000000000;
assign Upperletter[30] = 12'b111111111111;
assign Upperletter[31] = 12'b111111111111;
assign Upperletter[32] = 12'b111111111111;
assign Upperletter[33] = 12'b000000000000;
assign Upperletter[34] = 12'b111111111111;
assign Upperletter[35] = 12'b111111111111;
assign Upperletter[36] = 12'b111111111111;
assign Upperletter[37] = 12'b000000000000;
assign Upperletter[38] = 12'b111111111111;
assign Upperletter[39] = 12'b111111111111;
assign Upperletter[40] = 12'b111111111111;
assign Upperletter[41] = 12'b000000000000;
assign Upperletter[42] = 12'b111111111111;
assign Upperletter[43] = 12'b111111111111;
assign Upperletter[44] = 12'b111111111111;
assign Upperletter[45] = 12'b000000000000;
assign Upperletter[46] = 12'b111111111111;
assign Upperletter[47] = 12'b111111111111;
assign Upperletter[48] = 12'b111111111111;
assign Upperletter[49] = 12'b000000000000;
assign Upperletter[50] = 12'b111111111111;
assign Upperletter[51] = 12'b111111111111;
assign Upperletter[52] = 12'b111111111111;
assign Upperletter[53] = 12'b000000000000;
assign Upperletter[54] = 12'b111111111111;
assign Upperletter[55] = 12'b111111111111;
assign Upperletter[56] = 12'b111111111111;
assign Upperletter[57] = 12'b111111111111;
assign Upperletter[58] = 12'b111111111111;
assign Upperletter[59] = 12'b111111111111;
assign Upperletter[60] = 12'b111111111111;
assign Upperletter[61] = 12'b111111111111;
assign Upperletter[62] = 12'b111111111111;
assign Upperletter[63] = 12'b111111111111;
assign Upperletter[64] = 12'b111111111111;
assign Upperletter[65] = 12'b000000000000;
assign Upperletter[66] = 12'b000000000000;
assign Upperletter[67] = 12'b000000000000;
assign Upperletter[68] = 12'b000000000000;
assign Upperletter[69] = 12'b111111111111;
assign Upperletter[70] = 12'b111111111111;
assign Upperletter[71] = 12'b111111111111;
assign Upperletter[72] = 12'b111111111111;
assign Upperletter[73] = 12'b000000000000;
assign Upperletter[74] = 12'b111111111111;
assign Upperletter[75] = 12'b111111111111;
assign Upperletter[76] = 12'b111111111111;
assign Upperletter[77] = 12'b000000000000;
assign Upperletter[78] = 12'b111111111111;
assign Upperletter[79] = 12'b111111111111;
assign Upperletter[80] = 12'b111111111111;
assign Upperletter[81] = 12'b000000000000;
assign Upperletter[82] = 12'b111111111111;
assign Upperletter[83] = 12'b111111111111;
assign Upperletter[84] = 12'b111111111111;
assign Upperletter[85] = 12'b000000000000;
assign Upperletter[86] = 12'b111111111111;
assign Upperletter[87] = 12'b111111111111;
assign Upperletter[88] = 12'b111111111111;
assign Upperletter[89] = 12'b000000000000;
assign Upperletter[90] = 12'b000000000000;
assign Upperletter[91] = 12'b000000000000;
assign Upperletter[92] = 12'b000000000000;
assign Upperletter[93] = 12'b111111111111;
assign Upperletter[94] = 12'b111111111111;
assign Upperletter[95] = 12'b111111111111;
assign Upperletter[96] = 12'b111111111111;
assign Upperletter[97] = 12'b000000000000;
assign Upperletter[98] = 12'b111111111111;
assign Upperletter[99] = 12'b111111111111;
assign Upperletter[100] = 12'b111111111111;
assign Upperletter[101] = 12'b000000000000;
assign Upperletter[102] = 12'b111111111111;
assign Upperletter[103] = 12'b111111111111;
assign Upperletter[104] = 12'b111111111111;
assign Upperletter[105] = 12'b000000000000;
assign Upperletter[106] = 12'b111111111111;
assign Upperletter[107] = 12'b111111111111;
assign Upperletter[108] = 12'b111111111111;
assign Upperletter[109] = 12'b000000000000;
assign Upperletter[110] = 12'b111111111111;
assign Upperletter[111] = 12'b111111111111;
assign Upperletter[112] = 12'b111111111111;
assign Upperletter[113] = 12'b000000000000;
assign Upperletter[114] = 12'b000000000000;
assign Upperletter[115] = 12'b000000000000;
assign Upperletter[116] = 12'b000000000000;
assign Upperletter[117] = 12'b111111111111;
assign Upperletter[118] = 12'b111111111111;
assign Upperletter[119] = 12'b111111111111;
assign Upperletter[120] = 12'b111111111111;
assign Upperletter[121] = 12'b111111111111;
assign Upperletter[122] = 12'b111111111111;
assign Upperletter[123] = 12'b111111111111;
assign Upperletter[124] = 12'b111111111111;
assign Upperletter[125] = 12'b111111111111;
assign Upperletter[126] = 12'b111111111111;
assign Upperletter[127] = 12'b111111111111;
assign Upperletter[128] = 12'b111111111111;
assign Upperletter[129] = 12'b111111111111;
assign Upperletter[130] = 12'b000000000000;
assign Upperletter[131] = 12'b000000000000;
assign Upperletter[132] = 12'b000000000000;
assign Upperletter[133] = 12'b111111111111;
assign Upperletter[134] = 12'b111111111111;
assign Upperletter[135] = 12'b111111111111;
assign Upperletter[136] = 12'b111111111111;
assign Upperletter[137] = 12'b000000000000;
assign Upperletter[138] = 12'b111111111111;
assign Upperletter[139] = 12'b111111111111;
assign Upperletter[140] = 12'b111111111111;
assign Upperletter[141] = 12'b000000000000;
assign Upperletter[142] = 12'b111111111111;
assign Upperletter[143] = 12'b111111111111;
assign Upperletter[144] = 12'b111111111111;
assign Upperletter[145] = 12'b000000000000;
assign Upperletter[146] = 12'b111111111111;
assign Upperletter[147] = 12'b111111111111;
assign Upperletter[148] = 12'b111111111111;
assign Upperletter[149] = 12'b111111111111;
assign Upperletter[150] = 12'b111111111111;
assign Upperletter[151] = 12'b111111111111;
assign Upperletter[152] = 12'b111111111111;
assign Upperletter[153] = 12'b000000000000;
assign Upperletter[154] = 12'b111111111111;
assign Upperletter[155] = 12'b111111111111;
assign Upperletter[156] = 12'b111111111111;
assign Upperletter[157] = 12'b111111111111;
assign Upperletter[158] = 12'b111111111111;
assign Upperletter[159] = 12'b111111111111;
assign Upperletter[160] = 12'b111111111111;
assign Upperletter[161] = 12'b000000000000;
assign Upperletter[162] = 12'b111111111111;
assign Upperletter[163] = 12'b111111111111;
assign Upperletter[164] = 12'b111111111111;
assign Upperletter[165] = 12'b111111111111;
assign Upperletter[166] = 12'b111111111111;
assign Upperletter[167] = 12'b111111111111;
assign Upperletter[168] = 12'b111111111111;
assign Upperletter[169] = 12'b000000000000;
assign Upperletter[170] = 12'b111111111111;
assign Upperletter[171] = 12'b111111111111;
assign Upperletter[172] = 12'b111111111111;
assign Upperletter[173] = 12'b000000000000;
assign Upperletter[174] = 12'b111111111111;
assign Upperletter[175] = 12'b111111111111;
assign Upperletter[176] = 12'b111111111111;
assign Upperletter[177] = 12'b111111111111;
assign Upperletter[178] = 12'b000000000000;
assign Upperletter[179] = 12'b000000000000;
assign Upperletter[180] = 12'b000000000000;
assign Upperletter[181] = 12'b111111111111;
assign Upperletter[182] = 12'b111111111111;
assign Upperletter[183] = 12'b111111111111;
assign Upperletter[184] = 12'b111111111111;
assign Upperletter[185] = 12'b111111111111;
assign Upperletter[186] = 12'b111111111111;
assign Upperletter[187] = 12'b111111111111;
assign Upperletter[188] = 12'b111111111111;
assign Upperletter[189] = 12'b111111111111;
assign Upperletter[190] = 12'b111111111111;
assign Upperletter[191] = 12'b111111111111;
assign Upperletter[192] = 12'b111111111111;
assign Upperletter[193] = 12'b000000000000;
assign Upperletter[194] = 12'b000000000000;
assign Upperletter[195] = 12'b000000000000;
assign Upperletter[196] = 12'b000000000000;
assign Upperletter[197] = 12'b111111111111;
assign Upperletter[198] = 12'b111111111111;
assign Upperletter[199] = 12'b111111111111;
assign Upperletter[200] = 12'b111111111111;
assign Upperletter[201] = 12'b000000000000;
assign Upperletter[202] = 12'b111111111111;
assign Upperletter[203] = 12'b111111111111;
assign Upperletter[204] = 12'b111111111111;
assign Upperletter[205] = 12'b000000000000;
assign Upperletter[206] = 12'b111111111111;
assign Upperletter[207] = 12'b111111111111;
assign Upperletter[208] = 12'b111111111111;
assign Upperletter[209] = 12'b000000000000;
assign Upperletter[210] = 12'b111111111111;
assign Upperletter[211] = 12'b111111111111;
assign Upperletter[212] = 12'b111111111111;
assign Upperletter[213] = 12'b000000000000;
assign Upperletter[214] = 12'b111111111111;
assign Upperletter[215] = 12'b111111111111;
assign Upperletter[216] = 12'b111111111111;
assign Upperletter[217] = 12'b000000000000;
assign Upperletter[218] = 12'b111111111111;
assign Upperletter[219] = 12'b111111111111;
assign Upperletter[220] = 12'b111111111111;
assign Upperletter[221] = 12'b000000000000;
assign Upperletter[222] = 12'b111111111111;
assign Upperletter[223] = 12'b111111111111;
assign Upperletter[224] = 12'b111111111111;
assign Upperletter[225] = 12'b000000000000;
assign Upperletter[226] = 12'b111111111111;
assign Upperletter[227] = 12'b111111111111;
assign Upperletter[228] = 12'b111111111111;
assign Upperletter[229] = 12'b000000000000;
assign Upperletter[230] = 12'b111111111111;
assign Upperletter[231] = 12'b111111111111;
assign Upperletter[232] = 12'b111111111111;
assign Upperletter[233] = 12'b000000000000;
assign Upperletter[234] = 12'b111111111111;
assign Upperletter[235] = 12'b111111111111;
assign Upperletter[236] = 12'b111111111111;
assign Upperletter[237] = 12'b000000000000;
assign Upperletter[238] = 12'b111111111111;
assign Upperletter[239] = 12'b111111111111;
assign Upperletter[240] = 12'b111111111111;
assign Upperletter[241] = 12'b000000000000;
assign Upperletter[242] = 12'b000000000000;
assign Upperletter[243] = 12'b000000000000;
assign Upperletter[244] = 12'b000000000000;
assign Upperletter[245] = 12'b111111111111;
assign Upperletter[246] = 12'b111111111111;
assign Upperletter[247] = 12'b111111111111;
assign Upperletter[248] = 12'b111111111111;
assign Upperletter[249] = 12'b111111111111;
assign Upperletter[250] = 12'b111111111111;
assign Upperletter[251] = 12'b111111111111;
assign Upperletter[252] = 12'b111111111111;
assign Upperletter[253] = 12'b111111111111;
assign Upperletter[254] = 12'b111111111111;
assign Upperletter[255] = 12'b111111111111;
assign Upperletter[256] = 12'b111111111111;
assign Upperletter[257] = 12'b000000000000;
assign Upperletter[258] = 12'b000000000000;
assign Upperletter[259] = 12'b000000000000;
assign Upperletter[260] = 12'b000000000000;
assign Upperletter[261] = 12'b111111111111;
assign Upperletter[262] = 12'b111111111111;
assign Upperletter[263] = 12'b111111111111;
assign Upperletter[264] = 12'b111111111111;
assign Upperletter[265] = 12'b000000000000;
assign Upperletter[266] = 12'b111111111111;
assign Upperletter[267] = 12'b111111111111;
assign Upperletter[268] = 12'b111111111111;
assign Upperletter[269] = 12'b111111111111;
assign Upperletter[270] = 12'b111111111111;
assign Upperletter[271] = 12'b111111111111;
assign Upperletter[272] = 12'b111111111111;
assign Upperletter[273] = 12'b000000000000;
assign Upperletter[274] = 12'b111111111111;
assign Upperletter[275] = 12'b111111111111;
assign Upperletter[276] = 12'b111111111111;
assign Upperletter[277] = 12'b111111111111;
assign Upperletter[278] = 12'b111111111111;
assign Upperletter[279] = 12'b111111111111;
assign Upperletter[280] = 12'b111111111111;
assign Upperletter[281] = 12'b000000000000;
assign Upperletter[282] = 12'b000000000000;
assign Upperletter[283] = 12'b000000000000;
assign Upperletter[284] = 12'b111111111111;
assign Upperletter[285] = 12'b111111111111;
assign Upperletter[286] = 12'b111111111111;
assign Upperletter[287] = 12'b111111111111;
assign Upperletter[288] = 12'b111111111111;
assign Upperletter[289] = 12'b000000000000;
assign Upperletter[290] = 12'b111111111111;
assign Upperletter[291] = 12'b111111111111;
assign Upperletter[292] = 12'b111111111111;
assign Upperletter[293] = 12'b111111111111;
assign Upperletter[294] = 12'b111111111111;
assign Upperletter[295] = 12'b111111111111;
assign Upperletter[296] = 12'b111111111111;
assign Upperletter[297] = 12'b000000000000;
assign Upperletter[298] = 12'b111111111111;
assign Upperletter[299] = 12'b111111111111;
assign Upperletter[300] = 12'b111111111111;
assign Upperletter[301] = 12'b111111111111;
assign Upperletter[302] = 12'b111111111111;
assign Upperletter[303] = 12'b111111111111;
assign Upperletter[304] = 12'b111111111111;
assign Upperletter[305] = 12'b000000000000;
assign Upperletter[306] = 12'b000000000000;
assign Upperletter[307] = 12'b000000000000;
assign Upperletter[308] = 12'b000000000000;
assign Upperletter[309] = 12'b000000000000;
assign Upperletter[310] = 12'b111111111111;
assign Upperletter[311] = 12'b111111111111;
assign Upperletter[312] = 12'b111111111111;
assign Upperletter[313] = 12'b111111111111;
assign Upperletter[314] = 12'b111111111111;
assign Upperletter[315] = 12'b111111111111;
assign Upperletter[316] = 12'b111111111111;
assign Upperletter[317] = 12'b111111111111;
assign Upperletter[318] = 12'b111111111111;
assign Upperletter[319] = 12'b111111111111;
assign Upperletter[320] = 12'b111111111111;
assign Upperletter[321] = 12'b000000000000;
assign Upperletter[322] = 12'b000000000000;
assign Upperletter[323] = 12'b000000000000;
assign Upperletter[324] = 12'b000000000000;
assign Upperletter[325] = 12'b000000000000;
assign Upperletter[326] = 12'b111111111111;
assign Upperletter[327] = 12'b111111111111;
assign Upperletter[328] = 12'b111111111111;
assign Upperletter[329] = 12'b000000000000;
assign Upperletter[330] = 12'b111111111111;
assign Upperletter[331] = 12'b111111111111;
assign Upperletter[332] = 12'b111111111111;
assign Upperletter[333] = 12'b111111111111;
assign Upperletter[334] = 12'b111111111111;
assign Upperletter[335] = 12'b111111111111;
assign Upperletter[336] = 12'b111111111111;
assign Upperletter[337] = 12'b000000000000;
assign Upperletter[338] = 12'b111111111111;
assign Upperletter[339] = 12'b111111111111;
assign Upperletter[340] = 12'b111111111111;
assign Upperletter[341] = 12'b111111111111;
assign Upperletter[342] = 12'b111111111111;
assign Upperletter[343] = 12'b111111111111;
assign Upperletter[344] = 12'b111111111111;
assign Upperletter[345] = 12'b000000000000;
assign Upperletter[346] = 12'b000000000000;
assign Upperletter[347] = 12'b000000000000;
assign Upperletter[348] = 12'b000000000000;
assign Upperletter[349] = 12'b111111111111;
assign Upperletter[350] = 12'b111111111111;
assign Upperletter[351] = 12'b111111111111;
assign Upperletter[352] = 12'b111111111111;
assign Upperletter[353] = 12'b000000000000;
assign Upperletter[354] = 12'b111111111111;
assign Upperletter[355] = 12'b111111111111;
assign Upperletter[356] = 12'b111111111111;
assign Upperletter[357] = 12'b111111111111;
assign Upperletter[358] = 12'b111111111111;
assign Upperletter[359] = 12'b111111111111;
assign Upperletter[360] = 12'b111111111111;
assign Upperletter[361] = 12'b000000000000;
assign Upperletter[362] = 12'b111111111111;
assign Upperletter[363] = 12'b111111111111;
assign Upperletter[364] = 12'b111111111111;
assign Upperletter[365] = 12'b111111111111;
assign Upperletter[366] = 12'b111111111111;
assign Upperletter[367] = 12'b111111111111;
assign Upperletter[368] = 12'b111111111111;
assign Upperletter[369] = 12'b000000000000;
assign Upperletter[370] = 12'b111111111111;
assign Upperletter[371] = 12'b111111111111;
assign Upperletter[372] = 12'b111111111111;
assign Upperletter[373] = 12'b111111111111;
assign Upperletter[374] = 12'b111111111111;
assign Upperletter[375] = 12'b111111111111;
assign Upperletter[376] = 12'b111111111111;
assign Upperletter[377] = 12'b111111111111;
assign Upperletter[378] = 12'b111111111111;
assign Upperletter[379] = 12'b111111111111;
assign Upperletter[380] = 12'b111111111111;
assign Upperletter[381] = 12'b111111111111;
assign Upperletter[382] = 12'b111111111111;
assign Upperletter[383] = 12'b111111111111;
assign Upperletter[384] = 12'b111111111111;
assign Upperletter[385] = 12'b111111111111;
assign Upperletter[386] = 12'b000000000000;
assign Upperletter[387] = 12'b000000000000;
assign Upperletter[388] = 12'b000000000000;
assign Upperletter[389] = 12'b111111111111;
assign Upperletter[390] = 12'b111111111111;
assign Upperletter[391] = 12'b111111111111;
assign Upperletter[392] = 12'b111111111111;
assign Upperletter[393] = 12'b000000000000;
assign Upperletter[394] = 12'b111111111111;
assign Upperletter[395] = 12'b111111111111;
assign Upperletter[396] = 12'b111111111111;
assign Upperletter[397] = 12'b111111111111;
assign Upperletter[398] = 12'b111111111111;
assign Upperletter[399] = 12'b111111111111;
assign Upperletter[400] = 12'b111111111111;
assign Upperletter[401] = 12'b000000000000;
assign Upperletter[402] = 12'b111111111111;
assign Upperletter[403] = 12'b111111111111;
assign Upperletter[404] = 12'b111111111111;
assign Upperletter[405] = 12'b111111111111;
assign Upperletter[406] = 12'b111111111111;
assign Upperletter[407] = 12'b111111111111;
assign Upperletter[408] = 12'b111111111111;
assign Upperletter[409] = 12'b000000000000;
assign Upperletter[410] = 12'b111111111111;
assign Upperletter[411] = 12'b111111111111;
assign Upperletter[412] = 12'b000000000000;
assign Upperletter[413] = 12'b000000000000;
assign Upperletter[414] = 12'b111111111111;
assign Upperletter[415] = 12'b111111111111;
assign Upperletter[416] = 12'b111111111111;
assign Upperletter[417] = 12'b000000000000;
assign Upperletter[418] = 12'b111111111111;
assign Upperletter[419] = 12'b111111111111;
assign Upperletter[420] = 12'b111111111111;
assign Upperletter[421] = 12'b000000000000;
assign Upperletter[422] = 12'b111111111111;
assign Upperletter[423] = 12'b111111111111;
assign Upperletter[424] = 12'b111111111111;
assign Upperletter[425] = 12'b000000000000;
assign Upperletter[426] = 12'b111111111111;
assign Upperletter[427] = 12'b111111111111;
assign Upperletter[428] = 12'b111111111111;
assign Upperletter[429] = 12'b000000000000;
assign Upperletter[430] = 12'b111111111111;
assign Upperletter[431] = 12'b111111111111;
assign Upperletter[432] = 12'b111111111111;
assign Upperletter[433] = 12'b111111111111;
assign Upperletter[434] = 12'b000000000000;
assign Upperletter[435] = 12'b000000000000;
assign Upperletter[436] = 12'b000000000000;
assign Upperletter[437] = 12'b111111111111;
assign Upperletter[438] = 12'b111111111111;
assign Upperletter[439] = 12'b111111111111;
assign Upperletter[440] = 12'b111111111111;
assign Upperletter[441] = 12'b111111111111;
assign Upperletter[442] = 12'b111111111111;
assign Upperletter[443] = 12'b111111111111;
assign Upperletter[444] = 12'b111111111111;
assign Upperletter[445] = 12'b111111111111;
assign Upperletter[446] = 12'b111111111111;
assign Upperletter[447] = 12'b111111111111;
assign Upperletter[448] = 12'b111111111111;
assign Upperletter[449] = 12'b000000000000;
assign Upperletter[450] = 12'b111111111111;
assign Upperletter[451] = 12'b111111111111;
assign Upperletter[452] = 12'b111111111111;
assign Upperletter[453] = 12'b000000000000;
assign Upperletter[454] = 12'b111111111111;
assign Upperletter[455] = 12'b111111111111;
assign Upperletter[456] = 12'b111111111111;
assign Upperletter[457] = 12'b000000000000;
assign Upperletter[458] = 12'b111111111111;
assign Upperletter[459] = 12'b111111111111;
assign Upperletter[460] = 12'b111111111111;
assign Upperletter[461] = 12'b000000000000;
assign Upperletter[462] = 12'b111111111111;
assign Upperletter[463] = 12'b111111111111;
assign Upperletter[464] = 12'b111111111111;
assign Upperletter[465] = 12'b000000000000;
assign Upperletter[466] = 12'b111111111111;
assign Upperletter[467] = 12'b111111111111;
assign Upperletter[468] = 12'b111111111111;
assign Upperletter[469] = 12'b000000000000;
assign Upperletter[470] = 12'b111111111111;
assign Upperletter[471] = 12'b111111111111;
assign Upperletter[472] = 12'b111111111111;
assign Upperletter[473] = 12'b000000000000;
assign Upperletter[474] = 12'b000000000000;
assign Upperletter[475] = 12'b000000000000;
assign Upperletter[476] = 12'b000000000000;
assign Upperletter[477] = 12'b000000000000;
assign Upperletter[478] = 12'b111111111111;
assign Upperletter[479] = 12'b111111111111;
assign Upperletter[480] = 12'b111111111111;
assign Upperletter[481] = 12'b000000000000;
assign Upperletter[482] = 12'b111111111111;
assign Upperletter[483] = 12'b111111111111;
assign Upperletter[484] = 12'b111111111111;
assign Upperletter[485] = 12'b000000000000;
assign Upperletter[486] = 12'b111111111111;
assign Upperletter[487] = 12'b111111111111;
assign Upperletter[488] = 12'b111111111111;
assign Upperletter[489] = 12'b000000000000;
assign Upperletter[490] = 12'b111111111111;
assign Upperletter[491] = 12'b111111111111;
assign Upperletter[492] = 12'b111111111111;
assign Upperletter[493] = 12'b000000000000;
assign Upperletter[494] = 12'b111111111111;
assign Upperletter[495] = 12'b111111111111;
assign Upperletter[496] = 12'b111111111111;
assign Upperletter[497] = 12'b000000000000;
assign Upperletter[498] = 12'b111111111111;
assign Upperletter[499] = 12'b111111111111;
assign Upperletter[500] = 12'b111111111111;
assign Upperletter[501] = 12'b000000000000;
assign Upperletter[502] = 12'b111111111111;
assign Upperletter[503] = 12'b111111111111;
assign Upperletter[504] = 12'b111111111111;
assign Upperletter[505] = 12'b111111111111;
assign Upperletter[506] = 12'b111111111111;
assign Upperletter[507] = 12'b111111111111;
assign Upperletter[508] = 12'b111111111111;
assign Upperletter[509] = 12'b111111111111;
assign Upperletter[510] = 12'b111111111111;
assign Upperletter[511] = 12'b111111111111;
assign Upperletter[512] = 12'b111111111111;
assign Upperletter[513] = 12'b111111111111;
assign Upperletter[514] = 12'b000000000000;
assign Upperletter[515] = 12'b000000000000;
assign Upperletter[516] = 12'b000000000000;
assign Upperletter[517] = 12'b111111111111;
assign Upperletter[518] = 12'b111111111111;
assign Upperletter[519] = 12'b111111111111;
assign Upperletter[520] = 12'b111111111111;
assign Upperletter[521] = 12'b111111111111;
assign Upperletter[522] = 12'b111111111111;
assign Upperletter[523] = 12'b000000000000;
assign Upperletter[524] = 12'b111111111111;
assign Upperletter[525] = 12'b111111111111;
assign Upperletter[526] = 12'b111111111111;
assign Upperletter[527] = 12'b111111111111;
assign Upperletter[528] = 12'b111111111111;
assign Upperletter[529] = 12'b111111111111;
assign Upperletter[530] = 12'b111111111111;
assign Upperletter[531] = 12'b000000000000;
assign Upperletter[532] = 12'b111111111111;
assign Upperletter[533] = 12'b111111111111;
assign Upperletter[534] = 12'b111111111111;
assign Upperletter[535] = 12'b111111111111;
assign Upperletter[536] = 12'b111111111111;
assign Upperletter[537] = 12'b111111111111;
assign Upperletter[538] = 12'b111111111111;
assign Upperletter[539] = 12'b000000000000;
assign Upperletter[540] = 12'b111111111111;
assign Upperletter[541] = 12'b111111111111;
assign Upperletter[542] = 12'b111111111111;
assign Upperletter[543] = 12'b111111111111;
assign Upperletter[544] = 12'b111111111111;
assign Upperletter[545] = 12'b111111111111;
assign Upperletter[546] = 12'b111111111111;
assign Upperletter[547] = 12'b000000000000;
assign Upperletter[548] = 12'b111111111111;
assign Upperletter[549] = 12'b111111111111;
assign Upperletter[550] = 12'b111111111111;
assign Upperletter[551] = 12'b111111111111;
assign Upperletter[552] = 12'b111111111111;
assign Upperletter[553] = 12'b111111111111;
assign Upperletter[554] = 12'b111111111111;
assign Upperletter[555] = 12'b000000000000;
assign Upperletter[556] = 12'b111111111111;
assign Upperletter[557] = 12'b111111111111;
assign Upperletter[558] = 12'b111111111111;
assign Upperletter[559] = 12'b111111111111;
assign Upperletter[560] = 12'b111111111111;
assign Upperletter[561] = 12'b111111111111;
assign Upperletter[562] = 12'b000000000000;
assign Upperletter[563] = 12'b000000000000;
assign Upperletter[564] = 12'b000000000000;
assign Upperletter[565] = 12'b111111111111;
assign Upperletter[566] = 12'b111111111111;
assign Upperletter[567] = 12'b111111111111;
assign Upperletter[568] = 12'b111111111111;
assign Upperletter[569] = 12'b111111111111;
assign Upperletter[570] = 12'b111111111111;
assign Upperletter[571] = 12'b111111111111;
assign Upperletter[572] = 12'b111111111111;
assign Upperletter[573] = 12'b111111111111;
assign Upperletter[574] = 12'b111111111111;
assign Upperletter[575] = 12'b111111111111;
assign Upperletter[576] = 12'b111111111111;
assign Upperletter[577] = 12'b111111111111;
assign Upperletter[578] = 12'b111111111111;
assign Upperletter[579] = 12'b111111111111;
assign Upperletter[580] = 12'b000000000000;
assign Upperletter[581] = 12'b111111111111;
assign Upperletter[582] = 12'b111111111111;
assign Upperletter[583] = 12'b111111111111;
assign Upperletter[584] = 12'b111111111111;
assign Upperletter[585] = 12'b111111111111;
assign Upperletter[586] = 12'b111111111111;
assign Upperletter[587] = 12'b111111111111;
assign Upperletter[588] = 12'b000000000000;
assign Upperletter[589] = 12'b111111111111;
assign Upperletter[590] = 12'b111111111111;
assign Upperletter[591] = 12'b111111111111;
assign Upperletter[592] = 12'b111111111111;
assign Upperletter[593] = 12'b111111111111;
assign Upperletter[594] = 12'b111111111111;
assign Upperletter[595] = 12'b111111111111;
assign Upperletter[596] = 12'b000000000000;
assign Upperletter[597] = 12'b111111111111;
assign Upperletter[598] = 12'b111111111111;
assign Upperletter[599] = 12'b111111111111;
assign Upperletter[600] = 12'b111111111111;
assign Upperletter[601] = 12'b111111111111;
assign Upperletter[602] = 12'b111111111111;
assign Upperletter[603] = 12'b111111111111;
assign Upperletter[604] = 12'b000000000000;
assign Upperletter[605] = 12'b111111111111;
assign Upperletter[606] = 12'b111111111111;
assign Upperletter[607] = 12'b111111111111;
assign Upperletter[608] = 12'b111111111111;
assign Upperletter[609] = 12'b111111111111;
assign Upperletter[610] = 12'b111111111111;
assign Upperletter[611] = 12'b111111111111;
assign Upperletter[612] = 12'b000000000000;
assign Upperletter[613] = 12'b111111111111;
assign Upperletter[614] = 12'b111111111111;
assign Upperletter[615] = 12'b111111111111;
assign Upperletter[616] = 12'b111111111111;
assign Upperletter[617] = 12'b000000000000;
assign Upperletter[618] = 12'b111111111111;
assign Upperletter[619] = 12'b111111111111;
assign Upperletter[620] = 12'b000000000000;
assign Upperletter[621] = 12'b111111111111;
assign Upperletter[622] = 12'b111111111111;
assign Upperletter[623] = 12'b111111111111;
assign Upperletter[624] = 12'b111111111111;
assign Upperletter[625] = 12'b111111111111;
assign Upperletter[626] = 12'b000000000000;
assign Upperletter[627] = 12'b000000000000;
assign Upperletter[628] = 12'b111111111111;
assign Upperletter[629] = 12'b111111111111;
assign Upperletter[630] = 12'b111111111111;
assign Upperletter[631] = 12'b111111111111;
assign Upperletter[632] = 12'b111111111111;
assign Upperletter[633] = 12'b111111111111;
assign Upperletter[634] = 12'b111111111111;
assign Upperletter[635] = 12'b111111111111;
assign Upperletter[636] = 12'b111111111111;
assign Upperletter[637] = 12'b111111111111;
assign Upperletter[638] = 12'b111111111111;
assign Upperletter[639] = 12'b111111111111;
assign Upperletter[640] = 12'b111111111111;
assign Upperletter[641] = 12'b000000000000;
assign Upperletter[642] = 12'b111111111111;
assign Upperletter[643] = 12'b111111111111;
assign Upperletter[644] = 12'b111111111111;
assign Upperletter[645] = 12'b111111111111;
assign Upperletter[646] = 12'b111111111111;
assign Upperletter[647] = 12'b111111111111;
assign Upperletter[648] = 12'b111111111111;
assign Upperletter[649] = 12'b000000000000;
assign Upperletter[650] = 12'b111111111111;
assign Upperletter[651] = 12'b111111111111;
assign Upperletter[652] = 12'b111111111111;
assign Upperletter[653] = 12'b000000000000;
assign Upperletter[654] = 12'b111111111111;
assign Upperletter[655] = 12'b111111111111;
assign Upperletter[656] = 12'b111111111111;
assign Upperletter[657] = 12'b000000000000;
assign Upperletter[658] = 12'b111111111111;
assign Upperletter[659] = 12'b111111111111;
assign Upperletter[660] = 12'b000000000000;
assign Upperletter[661] = 12'b111111111111;
assign Upperletter[662] = 12'b111111111111;
assign Upperletter[663] = 12'b111111111111;
assign Upperletter[664] = 12'b111111111111;
assign Upperletter[665] = 12'b000000000000;
assign Upperletter[666] = 12'b000000000000;
assign Upperletter[667] = 12'b000000000000;
assign Upperletter[668] = 12'b111111111111;
assign Upperletter[669] = 12'b111111111111;
assign Upperletter[670] = 12'b111111111111;
assign Upperletter[671] = 12'b111111111111;
assign Upperletter[672] = 12'b111111111111;
assign Upperletter[673] = 12'b000000000000;
assign Upperletter[674] = 12'b111111111111;
assign Upperletter[675] = 12'b111111111111;
assign Upperletter[676] = 12'b000000000000;
assign Upperletter[677] = 12'b111111111111;
assign Upperletter[678] = 12'b111111111111;
assign Upperletter[679] = 12'b111111111111;
assign Upperletter[680] = 12'b111111111111;
assign Upperletter[681] = 12'b000000000000;
assign Upperletter[682] = 12'b111111111111;
assign Upperletter[683] = 12'b111111111111;
assign Upperletter[684] = 12'b111111111111;
assign Upperletter[685] = 12'b000000000000;
assign Upperletter[686] = 12'b111111111111;
assign Upperletter[687] = 12'b111111111111;
assign Upperletter[688] = 12'b111111111111;
assign Upperletter[689] = 12'b000000000000;
assign Upperletter[690] = 12'b111111111111;
assign Upperletter[691] = 12'b111111111111;
assign Upperletter[692] = 12'b111111111111;
assign Upperletter[693] = 12'b000000000000;
assign Upperletter[694] = 12'b111111111111;
assign Upperletter[695] = 12'b111111111111;
assign Upperletter[696] = 12'b111111111111;
assign Upperletter[697] = 12'b111111111111;
assign Upperletter[698] = 12'b111111111111;
assign Upperletter[699] = 12'b111111111111;
assign Upperletter[700] = 12'b111111111111;
assign Upperletter[701] = 12'b111111111111;
assign Upperletter[702] = 12'b111111111111;
assign Upperletter[703] = 12'b111111111111;
assign Upperletter[704] = 12'b111111111111;
assign Upperletter[705] = 12'b000000000000;
assign Upperletter[706] = 12'b111111111111;
assign Upperletter[707] = 12'b111111111111;
assign Upperletter[708] = 12'b111111111111;
assign Upperletter[709] = 12'b111111111111;
assign Upperletter[710] = 12'b111111111111;
assign Upperletter[711] = 12'b111111111111;
assign Upperletter[712] = 12'b111111111111;
assign Upperletter[713] = 12'b000000000000;
assign Upperletter[714] = 12'b111111111111;
assign Upperletter[715] = 12'b111111111111;
assign Upperletter[716] = 12'b111111111111;
assign Upperletter[717] = 12'b111111111111;
assign Upperletter[718] = 12'b111111111111;
assign Upperletter[719] = 12'b111111111111;
assign Upperletter[720] = 12'b111111111111;
assign Upperletter[721] = 12'b000000000000;
assign Upperletter[722] = 12'b111111111111;
assign Upperletter[723] = 12'b111111111111;
assign Upperletter[724] = 12'b111111111111;
assign Upperletter[725] = 12'b111111111111;
assign Upperletter[726] = 12'b111111111111;
assign Upperletter[727] = 12'b111111111111;
assign Upperletter[728] = 12'b111111111111;
assign Upperletter[729] = 12'b000000000000;
assign Upperletter[730] = 12'b111111111111;
assign Upperletter[731] = 12'b111111111111;
assign Upperletter[732] = 12'b111111111111;
assign Upperletter[733] = 12'b111111111111;
assign Upperletter[734] = 12'b111111111111;
assign Upperletter[735] = 12'b111111111111;
assign Upperletter[736] = 12'b111111111111;
assign Upperletter[737] = 12'b000000000000;
assign Upperletter[738] = 12'b111111111111;
assign Upperletter[739] = 12'b111111111111;
assign Upperletter[740] = 12'b111111111111;
assign Upperletter[741] = 12'b111111111111;
assign Upperletter[742] = 12'b111111111111;
assign Upperletter[743] = 12'b111111111111;
assign Upperletter[744] = 12'b111111111111;
assign Upperletter[745] = 12'b000000000000;
assign Upperletter[746] = 12'b111111111111;
assign Upperletter[747] = 12'b111111111111;
assign Upperletter[748] = 12'b111111111111;
assign Upperletter[749] = 12'b111111111111;
assign Upperletter[750] = 12'b111111111111;
assign Upperletter[751] = 12'b111111111111;
assign Upperletter[752] = 12'b111111111111;
assign Upperletter[753] = 12'b000000000000;
assign Upperletter[754] = 12'b000000000000;
assign Upperletter[755] = 12'b000000000000;
assign Upperletter[756] = 12'b000000000000;
assign Upperletter[757] = 12'b000000000000;
assign Upperletter[758] = 12'b111111111111;
assign Upperletter[759] = 12'b111111111111;
assign Upperletter[760] = 12'b111111111111;
assign Upperletter[761] = 12'b111111111111;
assign Upperletter[762] = 12'b111111111111;
assign Upperletter[763] = 12'b111111111111;
assign Upperletter[764] = 12'b111111111111;
assign Upperletter[765] = 12'b111111111111;
assign Upperletter[766] = 12'b111111111111;
assign Upperletter[767] = 12'b111111111111;
assign Upperletter[768] = 12'b111111111111;
assign Upperletter[769] = 12'b000000000000;
assign Upperletter[770] = 12'b111111111111;
assign Upperletter[771] = 12'b111111111111;
assign Upperletter[772] = 12'b111111111111;
assign Upperletter[773] = 12'b000000000000;
assign Upperletter[774] = 12'b111111111111;
assign Upperletter[775] = 12'b111111111111;
assign Upperletter[776] = 12'b111111111111;
assign Upperletter[777] = 12'b000000000000;
assign Upperletter[778] = 12'b000000000000;
assign Upperletter[779] = 12'b111111111111;
assign Upperletter[780] = 12'b000000000000;
assign Upperletter[781] = 12'b000000000000;
assign Upperletter[782] = 12'b111111111111;
assign Upperletter[783] = 12'b111111111111;
assign Upperletter[784] = 12'b111111111111;
assign Upperletter[785] = 12'b000000000000;
assign Upperletter[786] = 12'b111111111111;
assign Upperletter[787] = 12'b000000000000;
assign Upperletter[788] = 12'b111111111111;
assign Upperletter[789] = 12'b000000000000;
assign Upperletter[790] = 12'b111111111111;
assign Upperletter[791] = 12'b111111111111;
assign Upperletter[792] = 12'b111111111111;
assign Upperletter[793] = 12'b000000000000;
assign Upperletter[794] = 12'b111111111111;
assign Upperletter[795] = 12'b111111111111;
assign Upperletter[796] = 12'b111111111111;
assign Upperletter[797] = 12'b000000000000;
assign Upperletter[798] = 12'b111111111111;
assign Upperletter[799] = 12'b111111111111;
assign Upperletter[800] = 12'b111111111111;
assign Upperletter[801] = 12'b000000000000;
assign Upperletter[802] = 12'b111111111111;
assign Upperletter[803] = 12'b111111111111;
assign Upperletter[804] = 12'b111111111111;
assign Upperletter[805] = 12'b000000000000;
assign Upperletter[806] = 12'b111111111111;
assign Upperletter[807] = 12'b111111111111;
assign Upperletter[808] = 12'b111111111111;
assign Upperletter[809] = 12'b000000000000;
assign Upperletter[810] = 12'b111111111111;
assign Upperletter[811] = 12'b111111111111;
assign Upperletter[812] = 12'b111111111111;
assign Upperletter[813] = 12'b000000000000;
assign Upperletter[814] = 12'b111111111111;
assign Upperletter[815] = 12'b111111111111;
assign Upperletter[816] = 12'b111111111111;
assign Upperletter[817] = 12'b000000000000;
assign Upperletter[818] = 12'b111111111111;
assign Upperletter[819] = 12'b111111111111;
assign Upperletter[820] = 12'b111111111111;
assign Upperletter[821] = 12'b000000000000;
assign Upperletter[822] = 12'b111111111111;
assign Upperletter[823] = 12'b111111111111;
assign Upperletter[824] = 12'b111111111111;
assign Upperletter[825] = 12'b111111111111;
assign Upperletter[826] = 12'b111111111111;
assign Upperletter[827] = 12'b111111111111;
assign Upperletter[828] = 12'b111111111111;
assign Upperletter[829] = 12'b111111111111;
assign Upperletter[830] = 12'b111111111111;
assign Upperletter[831] = 12'b111111111111;
assign Upperletter[832] = 12'b111111111111;
assign Upperletter[833] = 12'b000000000000;
assign Upperletter[834] = 12'b111111111111;
assign Upperletter[835] = 12'b111111111111;
assign Upperletter[836] = 12'b111111111111;
assign Upperletter[837] = 12'b000000000000;
assign Upperletter[838] = 12'b111111111111;
assign Upperletter[839] = 12'b111111111111;
assign Upperletter[840] = 12'b111111111111;
assign Upperletter[841] = 12'b000000000000;
assign Upperletter[842] = 12'b000000000000;
assign Upperletter[843] = 12'b111111111111;
assign Upperletter[844] = 12'b111111111111;
assign Upperletter[845] = 12'b000000000000;
assign Upperletter[846] = 12'b111111111111;
assign Upperletter[847] = 12'b111111111111;
assign Upperletter[848] = 12'b111111111111;
assign Upperletter[849] = 12'b000000000000;
assign Upperletter[850] = 12'b111111111111;
assign Upperletter[851] = 12'b000000000000;
assign Upperletter[852] = 12'b111111111111;
assign Upperletter[853] = 12'b000000000000;
assign Upperletter[854] = 12'b111111111111;
assign Upperletter[855] = 12'b111111111111;
assign Upperletter[856] = 12'b111111111111;
assign Upperletter[857] = 12'b000000000000;
assign Upperletter[858] = 12'b111111111111;
assign Upperletter[859] = 12'b111111111111;
assign Upperletter[860] = 12'b000000000000;
assign Upperletter[861] = 12'b000000000000;
assign Upperletter[862] = 12'b111111111111;
assign Upperletter[863] = 12'b111111111111;
assign Upperletter[864] = 12'b111111111111;
assign Upperletter[865] = 12'b000000000000;
assign Upperletter[866] = 12'b111111111111;
assign Upperletter[867] = 12'b111111111111;
assign Upperletter[868] = 12'b111111111111;
assign Upperletter[869] = 12'b000000000000;
assign Upperletter[870] = 12'b111111111111;
assign Upperletter[871] = 12'b111111111111;
assign Upperletter[872] = 12'b111111111111;
assign Upperletter[873] = 12'b000000000000;
assign Upperletter[874] = 12'b111111111111;
assign Upperletter[875] = 12'b111111111111;
assign Upperletter[876] = 12'b111111111111;
assign Upperletter[877] = 12'b000000000000;
assign Upperletter[878] = 12'b111111111111;
assign Upperletter[879] = 12'b111111111111;
assign Upperletter[880] = 12'b111111111111;
assign Upperletter[881] = 12'b000000000000;
assign Upperletter[882] = 12'b111111111111;
assign Upperletter[883] = 12'b111111111111;
assign Upperletter[884] = 12'b111111111111;
assign Upperletter[885] = 12'b000000000000;
assign Upperletter[886] = 12'b111111111111;
assign Upperletter[887] = 12'b111111111111;
assign Upperletter[888] = 12'b111111111111;
assign Upperletter[889] = 12'b111111111111;
assign Upperletter[890] = 12'b111111111111;
assign Upperletter[891] = 12'b111111111111;
assign Upperletter[892] = 12'b111111111111;
assign Upperletter[893] = 12'b111111111111;
assign Upperletter[894] = 12'b111111111111;
assign Upperletter[895] = 12'b111111111111;
assign Upperletter[896] = 12'b111111111111;
assign Upperletter[897] = 12'b111111111111;
assign Upperletter[898] = 12'b000000000000;
assign Upperletter[899] = 12'b000000000000;
assign Upperletter[900] = 12'b000000000000;
assign Upperletter[901] = 12'b111111111111;
assign Upperletter[902] = 12'b111111111111;
assign Upperletter[903] = 12'b111111111111;
assign Upperletter[904] = 12'b111111111111;
assign Upperletter[905] = 12'b000000000000;
assign Upperletter[906] = 12'b111111111111;
assign Upperletter[907] = 12'b111111111111;
assign Upperletter[908] = 12'b111111111111;
assign Upperletter[909] = 12'b000000000000;
assign Upperletter[910] = 12'b111111111111;
assign Upperletter[911] = 12'b111111111111;
assign Upperletter[912] = 12'b111111111111;
assign Upperletter[913] = 12'b000000000000;
assign Upperletter[914] = 12'b111111111111;
assign Upperletter[915] = 12'b111111111111;
assign Upperletter[916] = 12'b111111111111;
assign Upperletter[917] = 12'b000000000000;
assign Upperletter[918] = 12'b111111111111;
assign Upperletter[919] = 12'b111111111111;
assign Upperletter[920] = 12'b111111111111;
assign Upperletter[921] = 12'b000000000000;
assign Upperletter[922] = 12'b111111111111;
assign Upperletter[923] = 12'b111111111111;
assign Upperletter[924] = 12'b111111111111;
assign Upperletter[925] = 12'b000000000000;
assign Upperletter[926] = 12'b111111111111;
assign Upperletter[927] = 12'b111111111111;
assign Upperletter[928] = 12'b111111111111;
assign Upperletter[929] = 12'b000000000000;
assign Upperletter[930] = 12'b111111111111;
assign Upperletter[931] = 12'b111111111111;
assign Upperletter[932] = 12'b111111111111;
assign Upperletter[933] = 12'b000000000000;
assign Upperletter[934] = 12'b111111111111;
assign Upperletter[935] = 12'b111111111111;
assign Upperletter[936] = 12'b111111111111;
assign Upperletter[937] = 12'b000000000000;
assign Upperletter[938] = 12'b111111111111;
assign Upperletter[939] = 12'b111111111111;
assign Upperletter[940] = 12'b111111111111;
assign Upperletter[941] = 12'b000000000000;
assign Upperletter[942] = 12'b111111111111;
assign Upperletter[943] = 12'b111111111111;
assign Upperletter[944] = 12'b111111111111;
assign Upperletter[945] = 12'b111111111111;
assign Upperletter[946] = 12'b000000000000;
assign Upperletter[947] = 12'b000000000000;
assign Upperletter[948] = 12'b000000000000;
assign Upperletter[949] = 12'b111111111111;
assign Upperletter[950] = 12'b111111111111;
assign Upperletter[951] = 12'b111111111111;
assign Upperletter[952] = 12'b111111111111;
assign Upperletter[953] = 12'b111111111111;
assign Upperletter[954] = 12'b111111111111;
assign Upperletter[955] = 12'b111111111111;
assign Upperletter[956] = 12'b111111111111;
assign Upperletter[957] = 12'b111111111111;
assign Upperletter[958] = 12'b111111111111;
assign Upperletter[959] = 12'b111111111111;
assign Upperletter[960] = 12'b111111111111;
assign Upperletter[961] = 12'b000000000000;
assign Upperletter[962] = 12'b000000000000;
assign Upperletter[963] = 12'b000000000000;
assign Upperletter[964] = 12'b000000000000;
assign Upperletter[965] = 12'b111111111111;
assign Upperletter[966] = 12'b111111111111;
assign Upperletter[967] = 12'b111111111111;
assign Upperletter[968] = 12'b111111111111;
assign Upperletter[969] = 12'b000000000000;
assign Upperletter[970] = 12'b111111111111;
assign Upperletter[971] = 12'b111111111111;
assign Upperletter[972] = 12'b111111111111;
assign Upperletter[973] = 12'b000000000000;
assign Upperletter[974] = 12'b111111111111;
assign Upperletter[975] = 12'b111111111111;
assign Upperletter[976] = 12'b111111111111;
assign Upperletter[977] = 12'b000000000000;
assign Upperletter[978] = 12'b111111111111;
assign Upperletter[979] = 12'b111111111111;
assign Upperletter[980] = 12'b111111111111;
assign Upperletter[981] = 12'b000000000000;
assign Upperletter[982] = 12'b111111111111;
assign Upperletter[983] = 12'b111111111111;
assign Upperletter[984] = 12'b111111111111;
assign Upperletter[985] = 12'b000000000000;
assign Upperletter[986] = 12'b000000000000;
assign Upperletter[987] = 12'b000000000000;
assign Upperletter[988] = 12'b000000000000;
assign Upperletter[989] = 12'b111111111111;
assign Upperletter[990] = 12'b111111111111;
assign Upperletter[991] = 12'b111111111111;
assign Upperletter[992] = 12'b111111111111;
assign Upperletter[993] = 12'b000000000000;
assign Upperletter[994] = 12'b111111111111;
assign Upperletter[995] = 12'b111111111111;
assign Upperletter[996] = 12'b111111111111;
assign Upperletter[997] = 12'b111111111111;
assign Upperletter[998] = 12'b111111111111;
assign Upperletter[999] = 12'b111111111111;
assign Upperletter[1000] = 12'b111111111111;
assign Upperletter[1001] = 12'b000000000000;
assign Upperletter[1002] = 12'b111111111111;
assign Upperletter[1003] = 12'b111111111111;
assign Upperletter[1004] = 12'b111111111111;
assign Upperletter[1005] = 12'b111111111111;
assign Upperletter[1006] = 12'b111111111111;
assign Upperletter[1007] = 12'b111111111111;
assign Upperletter[1008] = 12'b111111111111;
assign Upperletter[1009] = 12'b000000000000;
assign Upperletter[1010] = 12'b111111111111;
assign Upperletter[1011] = 12'b111111111111;
assign Upperletter[1012] = 12'b111111111111;
assign Upperletter[1013] = 12'b111111111111;
assign Upperletter[1014] = 12'b111111111111;
assign Upperletter[1015] = 12'b111111111111;
assign Upperletter[1016] = 12'b111111111111;
assign Upperletter[1017] = 12'b111111111111;
assign Upperletter[1018] = 12'b111111111111;
assign Upperletter[1019] = 12'b111111111111;
assign Upperletter[1020] = 12'b111111111111;
assign Upperletter[1021] = 12'b111111111111;
assign Upperletter[1022] = 12'b111111111111;
assign Upperletter[1023] = 12'b111111111111;
assign Upperletter[1024] = 12'b111111111111;
assign Upperletter[1025] = 12'b111111111111;
assign Upperletter[1026] = 12'b000000000000;
assign Upperletter[1027] = 12'b000000000000;
assign Upperletter[1028] = 12'b000000000000;
assign Upperletter[1029] = 12'b111111111111;
assign Upperletter[1030] = 12'b111111111111;
assign Upperletter[1031] = 12'b111111111111;
assign Upperletter[1032] = 12'b111111111111;
assign Upperletter[1033] = 12'b000000000000;
assign Upperletter[1034] = 12'b111111111111;
assign Upperletter[1035] = 12'b111111111111;
assign Upperletter[1036] = 12'b111111111111;
assign Upperletter[1037] = 12'b000000000000;
assign Upperletter[1038] = 12'b111111111111;
assign Upperletter[1039] = 12'b111111111111;
assign Upperletter[1040] = 12'b111111111111;
assign Upperletter[1041] = 12'b000000000000;
assign Upperletter[1042] = 12'b111111111111;
assign Upperletter[1043] = 12'b111111111111;
assign Upperletter[1044] = 12'b111111111111;
assign Upperletter[1045] = 12'b000000000000;
assign Upperletter[1046] = 12'b111111111111;
assign Upperletter[1047] = 12'b111111111111;
assign Upperletter[1048] = 12'b111111111111;
assign Upperletter[1049] = 12'b000000000000;
assign Upperletter[1050] = 12'b111111111111;
assign Upperletter[1051] = 12'b111111111111;
assign Upperletter[1052] = 12'b111111111111;
assign Upperletter[1053] = 12'b000000000000;
assign Upperletter[1054] = 12'b111111111111;
assign Upperletter[1055] = 12'b111111111111;
assign Upperletter[1056] = 12'b111111111111;
assign Upperletter[1057] = 12'b000000000000;
assign Upperletter[1058] = 12'b111111111111;
assign Upperletter[1059] = 12'b111111111111;
assign Upperletter[1060] = 12'b111111111111;
assign Upperletter[1061] = 12'b000000000000;
assign Upperletter[1062] = 12'b111111111111;
assign Upperletter[1063] = 12'b111111111111;
assign Upperletter[1064] = 12'b111111111111;
assign Upperletter[1065] = 12'b000000000000;
assign Upperletter[1066] = 12'b111111111111;
assign Upperletter[1067] = 12'b111111111111;
assign Upperletter[1068] = 12'b000000000000;
assign Upperletter[1069] = 12'b111111111111;
assign Upperletter[1070] = 12'b111111111111;
assign Upperletter[1071] = 12'b111111111111;
assign Upperletter[1072] = 12'b111111111111;
assign Upperletter[1073] = 12'b111111111111;
assign Upperletter[1074] = 12'b000000000000;
assign Upperletter[1075] = 12'b000000000000;
assign Upperletter[1076] = 12'b111111111111;
assign Upperletter[1077] = 12'b000000000000;
assign Upperletter[1078] = 12'b111111111111;
assign Upperletter[1079] = 12'b111111111111;
assign Upperletter[1080] = 12'b111111111111;
assign Upperletter[1081] = 12'b111111111111;
assign Upperletter[1082] = 12'b111111111111;
assign Upperletter[1083] = 12'b111111111111;
assign Upperletter[1084] = 12'b111111111111;
assign Upperletter[1085] = 12'b111111111111;
assign Upperletter[1086] = 12'b111111111111;
assign Upperletter[1087] = 12'b111111111111;
assign Upperletter[1088] = 12'b111111111111;
assign Upperletter[1089] = 12'b000000000000;
assign Upperletter[1090] = 12'b000000000000;
assign Upperletter[1091] = 12'b000000000000;
assign Upperletter[1092] = 12'b000000000000;
assign Upperletter[1093] = 12'b111111111111;
assign Upperletter[1094] = 12'b111111111111;
assign Upperletter[1095] = 12'b111111111111;
assign Upperletter[1096] = 12'b111111111111;
assign Upperletter[1097] = 12'b000000000000;
assign Upperletter[1098] = 12'b111111111111;
assign Upperletter[1099] = 12'b111111111111;
assign Upperletter[1100] = 12'b111111111111;
assign Upperletter[1101] = 12'b000000000000;
assign Upperletter[1102] = 12'b111111111111;
assign Upperletter[1103] = 12'b111111111111;
assign Upperletter[1104] = 12'b111111111111;
assign Upperletter[1105] = 12'b000000000000;
assign Upperletter[1106] = 12'b111111111111;
assign Upperletter[1107] = 12'b111111111111;
assign Upperletter[1108] = 12'b111111111111;
assign Upperletter[1109] = 12'b000000000000;
assign Upperletter[1110] = 12'b111111111111;
assign Upperletter[1111] = 12'b111111111111;
assign Upperletter[1112] = 12'b111111111111;
assign Upperletter[1113] = 12'b000000000000;
assign Upperletter[1114] = 12'b000000000000;
assign Upperletter[1115] = 12'b000000000000;
assign Upperletter[1116] = 12'b000000000000;
assign Upperletter[1117] = 12'b111111111111;
assign Upperletter[1118] = 12'b111111111111;
assign Upperletter[1119] = 12'b111111111111;
assign Upperletter[1120] = 12'b111111111111;
assign Upperletter[1121] = 12'b000000000000;
assign Upperletter[1122] = 12'b111111111111;
assign Upperletter[1123] = 12'b000000000000;
assign Upperletter[1124] = 12'b111111111111;
assign Upperletter[1125] = 12'b111111111111;
assign Upperletter[1126] = 12'b111111111111;
assign Upperletter[1127] = 12'b111111111111;
assign Upperletter[1128] = 12'b111111111111;
assign Upperletter[1129] = 12'b000000000000;
assign Upperletter[1130] = 12'b111111111111;
assign Upperletter[1131] = 12'b111111111111;
assign Upperletter[1132] = 12'b000000000000;
assign Upperletter[1133] = 12'b111111111111;
assign Upperletter[1134] = 12'b111111111111;
assign Upperletter[1135] = 12'b111111111111;
assign Upperletter[1136] = 12'b111111111111;
assign Upperletter[1137] = 12'b000000000000;
assign Upperletter[1138] = 12'b111111111111;
assign Upperletter[1139] = 12'b111111111111;
assign Upperletter[1140] = 12'b111111111111;
assign Upperletter[1141] = 12'b000000000000;
assign Upperletter[1142] = 12'b111111111111;
assign Upperletter[1143] = 12'b111111111111;
assign Upperletter[1144] = 12'b111111111111;
assign Upperletter[1145] = 12'b111111111111;
assign Upperletter[1146] = 12'b111111111111;
assign Upperletter[1147] = 12'b111111111111;
assign Upperletter[1148] = 12'b111111111111;
assign Upperletter[1149] = 12'b111111111111;
assign Upperletter[1150] = 12'b111111111111;
assign Upperletter[1151] = 12'b111111111111;
assign Upperletter[1152] = 12'b111111111111;
assign Upperletter[1153] = 12'b111111111111;
assign Upperletter[1154] = 12'b000000000000;
assign Upperletter[1155] = 12'b000000000000;
assign Upperletter[1156] = 12'b000000000000;
assign Upperletter[1157] = 12'b000000000000;
assign Upperletter[1158] = 12'b111111111111;
assign Upperletter[1159] = 12'b111111111111;
assign Upperletter[1160] = 12'b111111111111;
assign Upperletter[1161] = 12'b000000000000;
assign Upperletter[1162] = 12'b111111111111;
assign Upperletter[1163] = 12'b111111111111;
assign Upperletter[1164] = 12'b111111111111;
assign Upperletter[1165] = 12'b111111111111;
assign Upperletter[1166] = 12'b111111111111;
assign Upperletter[1167] = 12'b111111111111;
assign Upperletter[1168] = 12'b111111111111;
assign Upperletter[1169] = 12'b000000000000;
assign Upperletter[1170] = 12'b111111111111;
assign Upperletter[1171] = 12'b111111111111;
assign Upperletter[1172] = 12'b111111111111;
assign Upperletter[1173] = 12'b111111111111;
assign Upperletter[1174] = 12'b111111111111;
assign Upperletter[1175] = 12'b111111111111;
assign Upperletter[1176] = 12'b111111111111;
assign Upperletter[1177] = 12'b111111111111;
assign Upperletter[1178] = 12'b000000000000;
assign Upperletter[1179] = 12'b000000000000;
assign Upperletter[1180] = 12'b000000000000;
assign Upperletter[1181] = 12'b111111111111;
assign Upperletter[1182] = 12'b111111111111;
assign Upperletter[1183] = 12'b111111111111;
assign Upperletter[1184] = 12'b111111111111;
assign Upperletter[1185] = 12'b111111111111;
assign Upperletter[1186] = 12'b111111111111;
assign Upperletter[1187] = 12'b111111111111;
assign Upperletter[1188] = 12'b111111111111;
assign Upperletter[1189] = 12'b000000000000;
assign Upperletter[1190] = 12'b111111111111;
assign Upperletter[1191] = 12'b111111111111;
assign Upperletter[1192] = 12'b111111111111;
assign Upperletter[1193] = 12'b111111111111;
assign Upperletter[1194] = 12'b111111111111;
assign Upperletter[1195] = 12'b111111111111;
assign Upperletter[1196] = 12'b111111111111;
assign Upperletter[1197] = 12'b000000000000;
assign Upperletter[1198] = 12'b111111111111;
assign Upperletter[1199] = 12'b111111111111;
assign Upperletter[1200] = 12'b111111111111;
assign Upperletter[1201] = 12'b000000000000;
assign Upperletter[1202] = 12'b000000000000;
assign Upperletter[1203] = 12'b000000000000;
assign Upperletter[1204] = 12'b000000000000;
assign Upperletter[1205] = 12'b111111111111;
assign Upperletter[1206] = 12'b111111111111;
assign Upperletter[1207] = 12'b111111111111;
assign Upperletter[1208] = 12'b111111111111;
assign Upperletter[1209] = 12'b111111111111;
assign Upperletter[1210] = 12'b111111111111;
assign Upperletter[1211] = 12'b111111111111;
assign Upperletter[1212] = 12'b111111111111;
assign Upperletter[1213] = 12'b111111111111;
assign Upperletter[1214] = 12'b111111111111;
assign Upperletter[1215] = 12'b111111111111;
assign Upperletter[1216] = 12'b111111111111;
assign Upperletter[1217] = 12'b000000000000;
assign Upperletter[1218] = 12'b000000000000;
assign Upperletter[1219] = 12'b000000000000;
assign Upperletter[1220] = 12'b000000000000;
assign Upperletter[1221] = 12'b000000000000;
assign Upperletter[1222] = 12'b111111111111;
assign Upperletter[1223] = 12'b111111111111;
assign Upperletter[1224] = 12'b111111111111;
assign Upperletter[1225] = 12'b111111111111;
assign Upperletter[1226] = 12'b111111111111;
assign Upperletter[1227] = 12'b000000000000;
assign Upperletter[1228] = 12'b111111111111;
assign Upperletter[1229] = 12'b111111111111;
assign Upperletter[1230] = 12'b111111111111;
assign Upperletter[1231] = 12'b111111111111;
assign Upperletter[1232] = 12'b111111111111;
assign Upperletter[1233] = 12'b111111111111;
assign Upperletter[1234] = 12'b111111111111;
assign Upperletter[1235] = 12'b000000000000;
assign Upperletter[1236] = 12'b111111111111;
assign Upperletter[1237] = 12'b111111111111;
assign Upperletter[1238] = 12'b111111111111;
assign Upperletter[1239] = 12'b111111111111;
assign Upperletter[1240] = 12'b111111111111;
assign Upperletter[1241] = 12'b111111111111;
assign Upperletter[1242] = 12'b111111111111;
assign Upperletter[1243] = 12'b000000000000;
assign Upperletter[1244] = 12'b111111111111;
assign Upperletter[1245] = 12'b111111111111;
assign Upperletter[1246] = 12'b111111111111;
assign Upperletter[1247] = 12'b111111111111;
assign Upperletter[1248] = 12'b111111111111;
assign Upperletter[1249] = 12'b111111111111;
assign Upperletter[1250] = 12'b111111111111;
assign Upperletter[1251] = 12'b000000000000;
assign Upperletter[1252] = 12'b111111111111;
assign Upperletter[1253] = 12'b111111111111;
assign Upperletter[1254] = 12'b111111111111;
assign Upperletter[1255] = 12'b111111111111;
assign Upperletter[1256] = 12'b111111111111;
assign Upperletter[1257] = 12'b111111111111;
assign Upperletter[1258] = 12'b111111111111;
assign Upperletter[1259] = 12'b000000000000;
assign Upperletter[1260] = 12'b111111111111;
assign Upperletter[1261] = 12'b111111111111;
assign Upperletter[1262] = 12'b111111111111;
assign Upperletter[1263] = 12'b111111111111;
assign Upperletter[1264] = 12'b111111111111;
assign Upperletter[1265] = 12'b111111111111;
assign Upperletter[1266] = 12'b111111111111;
assign Upperletter[1267] = 12'b000000000000;
assign Upperletter[1268] = 12'b111111111111;
assign Upperletter[1269] = 12'b111111111111;
assign Upperletter[1270] = 12'b111111111111;
assign Upperletter[1271] = 12'b111111111111;
assign Upperletter[1272] = 12'b111111111111;
assign Upperletter[1273] = 12'b111111111111;
assign Upperletter[1274] = 12'b111111111111;
assign Upperletter[1275] = 12'b111111111111;
assign Upperletter[1276] = 12'b111111111111;
assign Upperletter[1277] = 12'b111111111111;
assign Upperletter[1278] = 12'b111111111111;
assign Upperletter[1279] = 12'b111111111111;
assign Upperletter[1280] = 12'b111111111111;
assign Upperletter[1281] = 12'b000000000000;
assign Upperletter[1282] = 12'b111111111111;
assign Upperletter[1283] = 12'b111111111111;
assign Upperletter[1284] = 12'b111111111111;
assign Upperletter[1285] = 12'b000000000000;
assign Upperletter[1286] = 12'b111111111111;
assign Upperletter[1287] = 12'b111111111111;
assign Upperletter[1288] = 12'b111111111111;
assign Upperletter[1289] = 12'b000000000000;
assign Upperletter[1290] = 12'b111111111111;
assign Upperletter[1291] = 12'b111111111111;
assign Upperletter[1292] = 12'b111111111111;
assign Upperletter[1293] = 12'b000000000000;
assign Upperletter[1294] = 12'b111111111111;
assign Upperletter[1295] = 12'b111111111111;
assign Upperletter[1296] = 12'b111111111111;
assign Upperletter[1297] = 12'b000000000000;
assign Upperletter[1298] = 12'b111111111111;
assign Upperletter[1299] = 12'b111111111111;
assign Upperletter[1300] = 12'b111111111111;
assign Upperletter[1301] = 12'b000000000000;
assign Upperletter[1302] = 12'b111111111111;
assign Upperletter[1303] = 12'b111111111111;
assign Upperletter[1304] = 12'b111111111111;
assign Upperletter[1305] = 12'b000000000000;
assign Upperletter[1306] = 12'b111111111111;
assign Upperletter[1307] = 12'b111111111111;
assign Upperletter[1308] = 12'b111111111111;
assign Upperletter[1309] = 12'b000000000000;
assign Upperletter[1310] = 12'b111111111111;
assign Upperletter[1311] = 12'b111111111111;
assign Upperletter[1312] = 12'b111111111111;
assign Upperletter[1313] = 12'b000000000000;
assign Upperletter[1314] = 12'b111111111111;
assign Upperletter[1315] = 12'b111111111111;
assign Upperletter[1316] = 12'b111111111111;
assign Upperletter[1317] = 12'b000000000000;
assign Upperletter[1318] = 12'b111111111111;
assign Upperletter[1319] = 12'b111111111111;
assign Upperletter[1320] = 12'b111111111111;
assign Upperletter[1321] = 12'b000000000000;
assign Upperletter[1322] = 12'b111111111111;
assign Upperletter[1323] = 12'b111111111111;
assign Upperletter[1324] = 12'b111111111111;
assign Upperletter[1325] = 12'b000000000000;
assign Upperletter[1326] = 12'b111111111111;
assign Upperletter[1327] = 12'b111111111111;
assign Upperletter[1328] = 12'b111111111111;
assign Upperletter[1329] = 12'b111111111111;
assign Upperletter[1330] = 12'b000000000000;
assign Upperletter[1331] = 12'b000000000000;
assign Upperletter[1332] = 12'b000000000000;
assign Upperletter[1333] = 12'b111111111111;
assign Upperletter[1334] = 12'b111111111111;
assign Upperletter[1335] = 12'b111111111111;
assign Upperletter[1336] = 12'b111111111111;
assign Upperletter[1337] = 12'b111111111111;
assign Upperletter[1338] = 12'b111111111111;
assign Upperletter[1339] = 12'b111111111111;
assign Upperletter[1340] = 12'b111111111111;
assign Upperletter[1341] = 12'b111111111111;
assign Upperletter[1342] = 12'b111111111111;
assign Upperletter[1343] = 12'b111111111111;
assign Upperletter[1344] = 12'b111111111111;
assign Upperletter[1345] = 12'b000000000000;
assign Upperletter[1346] = 12'b111111111111;
assign Upperletter[1347] = 12'b111111111111;
assign Upperletter[1348] = 12'b111111111111;
assign Upperletter[1349] = 12'b000000000000;
assign Upperletter[1350] = 12'b111111111111;
assign Upperletter[1351] = 12'b111111111111;
assign Upperletter[1352] = 12'b111111111111;
assign Upperletter[1353] = 12'b000000000000;
assign Upperletter[1354] = 12'b111111111111;
assign Upperletter[1355] = 12'b111111111111;
assign Upperletter[1356] = 12'b111111111111;
assign Upperletter[1357] = 12'b000000000000;
assign Upperletter[1358] = 12'b111111111111;
assign Upperletter[1359] = 12'b111111111111;
assign Upperletter[1360] = 12'b111111111111;
assign Upperletter[1361] = 12'b000000000000;
assign Upperletter[1362] = 12'b111111111111;
assign Upperletter[1363] = 12'b111111111111;
assign Upperletter[1364] = 12'b111111111111;
assign Upperletter[1365] = 12'b000000000000;
assign Upperletter[1366] = 12'b111111111111;
assign Upperletter[1367] = 12'b111111111111;
assign Upperletter[1368] = 12'b111111111111;
assign Upperletter[1369] = 12'b000000000000;
assign Upperletter[1370] = 12'b111111111111;
assign Upperletter[1371] = 12'b111111111111;
assign Upperletter[1372] = 12'b111111111111;
assign Upperletter[1373] = 12'b000000000000;
assign Upperletter[1374] = 12'b111111111111;
assign Upperletter[1375] = 12'b111111111111;
assign Upperletter[1376] = 12'b111111111111;
assign Upperletter[1377] = 12'b000000000000;
assign Upperletter[1378] = 12'b111111111111;
assign Upperletter[1379] = 12'b111111111111;
assign Upperletter[1380] = 12'b111111111111;
assign Upperletter[1381] = 12'b000000000000;
assign Upperletter[1382] = 12'b111111111111;
assign Upperletter[1383] = 12'b111111111111;
assign Upperletter[1384] = 12'b111111111111;
assign Upperletter[1385] = 12'b111111111111;
assign Upperletter[1386] = 12'b000000000000;
assign Upperletter[1387] = 12'b111111111111;
assign Upperletter[1388] = 12'b000000000000;
assign Upperletter[1389] = 12'b111111111111;
assign Upperletter[1390] = 12'b111111111111;
assign Upperletter[1391] = 12'b111111111111;
assign Upperletter[1392] = 12'b111111111111;
assign Upperletter[1393] = 12'b111111111111;
assign Upperletter[1394] = 12'b111111111111;
assign Upperletter[1395] = 12'b000000000000;
assign Upperletter[1396] = 12'b111111111111;
assign Upperletter[1397] = 12'b111111111111;
assign Upperletter[1398] = 12'b111111111111;
assign Upperletter[1399] = 12'b111111111111;
assign Upperletter[1400] = 12'b111111111111;
assign Upperletter[1401] = 12'b111111111111;
assign Upperletter[1402] = 12'b111111111111;
assign Upperletter[1403] = 12'b111111111111;
assign Upperletter[1404] = 12'b111111111111;
assign Upperletter[1405] = 12'b111111111111;
assign Upperletter[1406] = 12'b111111111111;
assign Upperletter[1407] = 12'b111111111111;
assign Upperletter[1408] = 12'b111111111111;
assign Upperletter[1409] = 12'b000000000000;
assign Upperletter[1410] = 12'b111111111111;
assign Upperletter[1411] = 12'b111111111111;
assign Upperletter[1412] = 12'b111111111111;
assign Upperletter[1413] = 12'b000000000000;
assign Upperletter[1414] = 12'b111111111111;
assign Upperletter[1415] = 12'b111111111111;
assign Upperletter[1416] = 12'b111111111111;
assign Upperletter[1417] = 12'b000000000000;
assign Upperletter[1418] = 12'b111111111111;
assign Upperletter[1419] = 12'b111111111111;
assign Upperletter[1420] = 12'b111111111111;
assign Upperletter[1421] = 12'b000000000000;
assign Upperletter[1422] = 12'b111111111111;
assign Upperletter[1423] = 12'b111111111111;
assign Upperletter[1424] = 12'b111111111111;
assign Upperletter[1425] = 12'b000000000000;
assign Upperletter[1426] = 12'b111111111111;
assign Upperletter[1427] = 12'b111111111111;
assign Upperletter[1428] = 12'b111111111111;
assign Upperletter[1429] = 12'b000000000000;
assign Upperletter[1430] = 12'b111111111111;
assign Upperletter[1431] = 12'b111111111111;
assign Upperletter[1432] = 12'b111111111111;
assign Upperletter[1433] = 12'b000000000000;
assign Upperletter[1434] = 12'b111111111111;
assign Upperletter[1435] = 12'b111111111111;
assign Upperletter[1436] = 12'b111111111111;
assign Upperletter[1437] = 12'b000000000000;
assign Upperletter[1438] = 12'b111111111111;
assign Upperletter[1439] = 12'b111111111111;
assign Upperletter[1440] = 12'b111111111111;
assign Upperletter[1441] = 12'b000000000000;
assign Upperletter[1442] = 12'b111111111111;
assign Upperletter[1443] = 12'b000000000000;
assign Upperletter[1444] = 12'b111111111111;
assign Upperletter[1445] = 12'b000000000000;
assign Upperletter[1446] = 12'b111111111111;
assign Upperletter[1447] = 12'b111111111111;
assign Upperletter[1448] = 12'b111111111111;
assign Upperletter[1449] = 12'b000000000000;
assign Upperletter[1450] = 12'b000000000000;
assign Upperletter[1451] = 12'b111111111111;
assign Upperletter[1452] = 12'b000000000000;
assign Upperletter[1453] = 12'b000000000000;
assign Upperletter[1454] = 12'b111111111111;
assign Upperletter[1455] = 12'b111111111111;
assign Upperletter[1456] = 12'b111111111111;
assign Upperletter[1457] = 12'b000000000000;
assign Upperletter[1458] = 12'b111111111111;
assign Upperletter[1459] = 12'b111111111111;
assign Upperletter[1460] = 12'b111111111111;
assign Upperletter[1461] = 12'b000000000000;
assign Upperletter[1462] = 12'b111111111111;
assign Upperletter[1463] = 12'b111111111111;
assign Upperletter[1464] = 12'b111111111111;
assign Upperletter[1465] = 12'b111111111111;
assign Upperletter[1466] = 12'b111111111111;
assign Upperletter[1467] = 12'b111111111111;
assign Upperletter[1468] = 12'b111111111111;
assign Upperletter[1469] = 12'b111111111111;
assign Upperletter[1470] = 12'b111111111111;
assign Upperletter[1471] = 12'b111111111111;
assign Upperletter[1472] = 12'b111111111111;
assign Upperletter[1473] = 12'b000000000000;
assign Upperletter[1474] = 12'b111111111111;
assign Upperletter[1475] = 12'b111111111111;
assign Upperletter[1476] = 12'b111111111111;
assign Upperletter[1477] = 12'b000000000000;
assign Upperletter[1478] = 12'b111111111111;
assign Upperletter[1479] = 12'b111111111111;
assign Upperletter[1480] = 12'b111111111111;
assign Upperletter[1481] = 12'b000000000000;
assign Upperletter[1482] = 12'b111111111111;
assign Upperletter[1483] = 12'b111111111111;
assign Upperletter[1484] = 12'b111111111111;
assign Upperletter[1485] = 12'b000000000000;
assign Upperletter[1486] = 12'b111111111111;
assign Upperletter[1487] = 12'b111111111111;
assign Upperletter[1488] = 12'b111111111111;
assign Upperletter[1489] = 12'b111111111111;
assign Upperletter[1490] = 12'b000000000000;
assign Upperletter[1491] = 12'b111111111111;
assign Upperletter[1492] = 12'b000000000000;
assign Upperletter[1493] = 12'b111111111111;
assign Upperletter[1494] = 12'b111111111111;
assign Upperletter[1495] = 12'b111111111111;
assign Upperletter[1496] = 12'b111111111111;
assign Upperletter[1497] = 12'b111111111111;
assign Upperletter[1498] = 12'b111111111111;
assign Upperletter[1499] = 12'b000000000000;
assign Upperletter[1500] = 12'b111111111111;
assign Upperletter[1501] = 12'b111111111111;
assign Upperletter[1502] = 12'b111111111111;
assign Upperletter[1503] = 12'b111111111111;
assign Upperletter[1504] = 12'b111111111111;
assign Upperletter[1505] = 12'b111111111111;
assign Upperletter[1506] = 12'b000000000000;
assign Upperletter[1507] = 12'b111111111111;
assign Upperletter[1508] = 12'b000000000000;
assign Upperletter[1509] = 12'b111111111111;
assign Upperletter[1510] = 12'b111111111111;
assign Upperletter[1511] = 12'b111111111111;
assign Upperletter[1512] = 12'b111111111111;
assign Upperletter[1513] = 12'b000000000000;
assign Upperletter[1514] = 12'b111111111111;
assign Upperletter[1515] = 12'b111111111111;
assign Upperletter[1516] = 12'b111111111111;
assign Upperletter[1517] = 12'b000000000000;
assign Upperletter[1518] = 12'b111111111111;
assign Upperletter[1519] = 12'b111111111111;
assign Upperletter[1520] = 12'b111111111111;
assign Upperletter[1521] = 12'b000000000000;
assign Upperletter[1522] = 12'b111111111111;
assign Upperletter[1523] = 12'b111111111111;
assign Upperletter[1524] = 12'b111111111111;
assign Upperletter[1525] = 12'b000000000000;
assign Upperletter[1526] = 12'b111111111111;
assign Upperletter[1527] = 12'b111111111111;
assign Upperletter[1528] = 12'b111111111111;
assign Upperletter[1529] = 12'b111111111111;
assign Upperletter[1530] = 12'b111111111111;
assign Upperletter[1531] = 12'b111111111111;
assign Upperletter[1532] = 12'b111111111111;
assign Upperletter[1533] = 12'b111111111111;
assign Upperletter[1534] = 12'b111111111111;
assign Upperletter[1535] = 12'b111111111111;
assign Upperletter[1536] = 12'b111111111111;
assign Upperletter[1537] = 12'b000000000000;
assign Upperletter[1538] = 12'b111111111111;
assign Upperletter[1539] = 12'b111111111111;
assign Upperletter[1540] = 12'b111111111111;
assign Upperletter[1541] = 12'b000000000000;
assign Upperletter[1542] = 12'b111111111111;
assign Upperletter[1543] = 12'b111111111111;
assign Upperletter[1544] = 12'b111111111111;
assign Upperletter[1545] = 12'b000000000000;
assign Upperletter[1546] = 12'b111111111111;
assign Upperletter[1547] = 12'b111111111111;
assign Upperletter[1548] = 12'b111111111111;
assign Upperletter[1549] = 12'b000000000000;
assign Upperletter[1550] = 12'b111111111111;
assign Upperletter[1551] = 12'b111111111111;
assign Upperletter[1552] = 12'b111111111111;
assign Upperletter[1553] = 12'b111111111111;
assign Upperletter[1554] = 12'b000000000000;
assign Upperletter[1555] = 12'b111111111111;
assign Upperletter[1556] = 12'b000000000000;
assign Upperletter[1557] = 12'b111111111111;
assign Upperletter[1558] = 12'b111111111111;
assign Upperletter[1559] = 12'b111111111111;
assign Upperletter[1560] = 12'b111111111111;
assign Upperletter[1561] = 12'b111111111111;
assign Upperletter[1562] = 12'b111111111111;
assign Upperletter[1563] = 12'b000000000000;
assign Upperletter[1564] = 12'b111111111111;
assign Upperletter[1565] = 12'b111111111111;
assign Upperletter[1566] = 12'b111111111111;
assign Upperletter[1567] = 12'b111111111111;
assign Upperletter[1568] = 12'b111111111111;
assign Upperletter[1569] = 12'b111111111111;
assign Upperletter[1570] = 12'b111111111111;
assign Upperletter[1571] = 12'b000000000000;
assign Upperletter[1572] = 12'b111111111111;
assign Upperletter[1573] = 12'b111111111111;
assign Upperletter[1574] = 12'b111111111111;
assign Upperletter[1575] = 12'b111111111111;
assign Upperletter[1576] = 12'b111111111111;
assign Upperletter[1577] = 12'b111111111111;
assign Upperletter[1578] = 12'b111111111111;
assign Upperletter[1579] = 12'b000000000000;
assign Upperletter[1580] = 12'b111111111111;
assign Upperletter[1581] = 12'b111111111111;
assign Upperletter[1582] = 12'b111111111111;
assign Upperletter[1583] = 12'b111111111111;
assign Upperletter[1584] = 12'b111111111111;
assign Upperletter[1585] = 12'b111111111111;
assign Upperletter[1586] = 12'b111111111111;
assign Upperletter[1587] = 12'b000000000000;
assign Upperletter[1588] = 12'b111111111111;
assign Upperletter[1589] = 12'b111111111111;
assign Upperletter[1590] = 12'b111111111111;
assign Upperletter[1591] = 12'b111111111111;
assign Upperletter[1592] = 12'b111111111111;
assign Upperletter[1593] = 12'b111111111111;
assign Upperletter[1594] = 12'b111111111111;
assign Upperletter[1595] = 12'b111111111111;
assign Upperletter[1596] = 12'b111111111111;
assign Upperletter[1597] = 12'b111111111111;
assign Upperletter[1598] = 12'b111111111111;
assign Upperletter[1599] = 12'b111111111111;
assign Upperletter[1600] = 12'b111111111111;
assign Upperletter[1601] = 12'b000000000000;
assign Upperletter[1602] = 12'b000000000000;
assign Upperletter[1603] = 12'b000000000000;
assign Upperletter[1604] = 12'b000000000000;
assign Upperletter[1605] = 12'b000000000000;
assign Upperletter[1606] = 12'b111111111111;
assign Upperletter[1607] = 12'b111111111111;
assign Upperletter[1608] = 12'b111111111111;
assign Upperletter[1609] = 12'b111111111111;
assign Upperletter[1610] = 12'b111111111111;
assign Upperletter[1611] = 12'b111111111111;
assign Upperletter[1612] = 12'b111111111111;
assign Upperletter[1613] = 12'b000000000000;
assign Upperletter[1614] = 12'b111111111111;
assign Upperletter[1615] = 12'b111111111111;
assign Upperletter[1616] = 12'b111111111111;
assign Upperletter[1617] = 12'b111111111111;
assign Upperletter[1618] = 12'b111111111111;
assign Upperletter[1619] = 12'b111111111111;
assign Upperletter[1620] = 12'b000000000000;
assign Upperletter[1621] = 12'b111111111111;
assign Upperletter[1622] = 12'b111111111111;
assign Upperletter[1623] = 12'b111111111111;
assign Upperletter[1624] = 12'b111111111111;
assign Upperletter[1625] = 12'b111111111111;
assign Upperletter[1626] = 12'b111111111111;
assign Upperletter[1627] = 12'b000000000000;
assign Upperletter[1628] = 12'b111111111111;
assign Upperletter[1629] = 12'b111111111111;
assign Upperletter[1630] = 12'b111111111111;
assign Upperletter[1631] = 12'b111111111111;
assign Upperletter[1632] = 12'b111111111111;
assign Upperletter[1633] = 12'b111111111111;
assign Upperletter[1634] = 12'b000000000000;
assign Upperletter[1635] = 12'b111111111111;
assign Upperletter[1636] = 12'b111111111111;
assign Upperletter[1637] = 12'b111111111111;
assign Upperletter[1638] = 12'b111111111111;
assign Upperletter[1639] = 12'b111111111111;
assign Upperletter[1640] = 12'b111111111111;
assign Upperletter[1641] = 12'b000000000000;
assign Upperletter[1642] = 12'b111111111111;
assign Upperletter[1643] = 12'b111111111111;
assign Upperletter[1644] = 12'b111111111111;
assign Upperletter[1645] = 12'b111111111111;
assign Upperletter[1646] = 12'b111111111111;
assign Upperletter[1647] = 12'b111111111111;
assign Upperletter[1648] = 12'b111111111111;
assign Upperletter[1649] = 12'b000000000000;
assign Upperletter[1650] = 12'b000000000000;
assign Upperletter[1651] = 12'b000000000000;
assign Upperletter[1652] = 12'b000000000000;
assign Upperletter[1653] = 12'b000000000000;
assign Upperletter[1654] = 12'b111111111111;
assign Upperletter[1655] = 12'b111111111111;
assign Upperletter[1656] = 12'b111111111111;
assign Upperletter[1657] = 12'b111111111111;
assign Upperletter[1658] = 12'b111111111111;
assign Upperletter[1659] = 12'b111111111111;
assign Upperletter[1660] = 12'b111111111111;
assign Upperletter[1661] = 12'b111111111111;
assign Upperletter[1662] = 12'b111111111111;
assign Upperletter[1663] = 12'b111111111111;
   
   
endmodule
