`timescale 1ns/1ps

module Decode_And_Exectue_t;
